library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity dadda is
	port (
		pp0: in std_logic_vector(63 downto 0);
		pp1: in std_logic_vector(63 downto 0);
		pp2: in std_logic_vector(63 downto 0);
		pp3: in std_logic_vector(63 downto 0);
		pp4: in std_logic_vector(63 downto 0);
		pp5: in std_logic_vector(63 downto 0);
		pp6: in std_logic_vector(63 downto 0);
		pp7: in std_logic_vector(63 downto 0);
		pp8: in std_logic_vector(63 downto 0);
		pp9: in std_logic_vector(63 downto 0);
		pp10: in std_logic_vector(63 downto 0);
		pp11: in std_logic_vector(63 downto 0);
		pp12: in std_logic_vector(63 downto 0);
		pp13: in std_logic_vector(63 downto 0);
		pp14: in std_logic_vector(63 downto 0);
		pp15: in std_logic_vector(63 downto 0);
		pp16: in std_logic_vector(63 downto 0);
		res: out std_logic_vector(63 downto 0)
	);
end entity dadda;

architecture structural of dadda is
	component ha is
		port (
			a: in std_logic;
			b: in std_logic;
			s: out std_logic;
			co: out std_logic
		);
	end component ha;

	component fa is
		port (
			a: in std_logic;
			b: in std_logic;
			ci: in std_logic;
			s: out std_logic;
			co: out std_logic
		);
	end component fa;

	type dadda6_arr is array(0 to 16) of std_logic_vector(63 downto 0);
	type dadda5_arr is array(0 to 12) of std_logic_vector(63 downto 0);
	type dadda4_arr is array(0 to 8) of std_logic_vector(63 downto 0);
	type dadda3_arr is array(0 to 5) of std_logic_vector(63 downto 0);
	type dadda2_arr is array(0 to 3) of std_logic_vector(63 downto 0);
	type dadda1_arr is array(0 to 2) of std_logic_vector(63 downto 0);
	type dadda0_arr is array(0 to 1) of std_logic_vector(63 downto 0);

	signal dadda_tree_6: dadda6_arr;
	signal dadda_tree_5: dadda5_arr;
	signal dadda_tree_4: dadda4_arr;
	signal dadda_tree_3: dadda3_arr;
	signal dadda_tree_2: dadda2_arr;
	signal dadda_tree_1: dadda1_arr;
	signal dadda_tree_0: dadda0_arr;

	signal res_ext: std_logic_vector(64 downto 0);
begin
	dadda_tree_6(0) <= pp0;
	dadda_tree_6(1) <= pp1;
	dadda_tree_6(2) <= pp2;
	dadda_tree_6(3) <= pp3;
	dadda_tree_6(4) <= pp4;
	dadda_tree_6(5) <= pp5;
	dadda_tree_6(6) <= pp6;
	dadda_tree_6(7) <= pp7;
	dadda_tree_6(8) <= pp8;
	dadda_tree_6(9) <= pp9;
	dadda_tree_6(10) <= pp10;
	dadda_tree_6(11) <= pp11;
	dadda_tree_6(12) <= pp12;
	dadda_tree_6(13) <= pp13;
	dadda_tree_6(14) <= pp14;
	dadda_tree_6(15) <= pp15;
	dadda_tree_6(16) <= pp16;

	res_ext <= std_logic_vector(unsigned(dadda_tree_0(0)) + unsigned(dadda_tree_0(1)))
	res <= res_ext(63 downto 0);

	

	-- AUTO-GENERATED CODE



	dadda_tree_5(0)(0) <= dadda_tree_6(0)(0);
	dadda_tree_5(1)(0) <= dadda_tree_6(1)(0);
	dadda_tree_5(0)(1) <= dadda_tree_6(0)(1);
	dadda_tree_5(0)(2) <= dadda_tree_6(0)(2);
	dadda_tree_5(1)(2) <= dadda_tree_6(1)(2);
	dadda_tree_5(2)(2) <= dadda_tree_6(2)(2);
	dadda_tree_5(0)(3) <= dadda_tree_6(0)(3);
	dadda_tree_5(1)(3) <= dadda_tree_6(1)(3);
	dadda_tree_5(0)(4) <= dadda_tree_6(0)(4);
	dadda_tree_5(1)(4) <= dadda_tree_6(1)(4);
	dadda_tree_5(2)(4) <= dadda_tree_6(2)(4);
	dadda_tree_5(3)(4) <= dadda_tree_6(3)(4);
	dadda_tree_5(0)(5) <= dadda_tree_6(0)(5);
	dadda_tree_5(1)(5) <= dadda_tree_6(1)(5);
	dadda_tree_5(2)(5) <= dadda_tree_6(2)(5);
	dadda_tree_5(0)(6) <= dadda_tree_6(0)(6);
	dadda_tree_5(1)(6) <= dadda_tree_6(1)(6);
	dadda_tree_5(2)(6) <= dadda_tree_6(2)(6);
	dadda_tree_5(3)(6) <= dadda_tree_6(3)(6);
	dadda_tree_5(4)(6) <= dadda_tree_6(4)(6);
	dadda_tree_5(0)(7) <= dadda_tree_6(0)(7);
	dadda_tree_5(1)(7) <= dadda_tree_6(1)(7);
	dadda_tree_5(2)(7) <= dadda_tree_6(2)(7);
	dadda_tree_5(3)(7) <= dadda_tree_6(3)(7);
	dadda_tree_5(0)(8) <= dadda_tree_6(0)(8);
	dadda_tree_5(1)(8) <= dadda_tree_6(1)(8);
	dadda_tree_5(2)(8) <= dadda_tree_6(2)(8);
	dadda_tree_5(3)(8) <= dadda_tree_6(3)(8);
	dadda_tree_5(4)(8) <= dadda_tree_6(4)(8);
	dadda_tree_5(5)(8) <= dadda_tree_6(5)(8);
	dadda_tree_5(0)(9) <= dadda_tree_6(0)(9);
	dadda_tree_5(1)(9) <= dadda_tree_6(1)(9);
	dadda_tree_5(2)(9) <= dadda_tree_6(2)(9);
	dadda_tree_5(3)(9) <= dadda_tree_6(3)(9);
	dadda_tree_5(4)(9) <= dadda_tree_6(4)(9);
	dadda_tree_5(0)(10) <= dadda_tree_6(0)(10);
	dadda_tree_5(1)(10) <= dadda_tree_6(1)(10);
	dadda_tree_5(2)(10) <= dadda_tree_6(2)(10);
	dadda_tree_5(3)(10) <= dadda_tree_6(3)(10);
	dadda_tree_5(4)(10) <= dadda_tree_6(4)(10);
	dadda_tree_5(5)(10) <= dadda_tree_6(5)(10);
	dadda_tree_5(6)(10) <= dadda_tree_6(6)(10);
	dadda_tree_5(0)(11) <= dadda_tree_6(0)(11);
	dadda_tree_5(1)(11) <= dadda_tree_6(1)(11);
	dadda_tree_5(2)(11) <= dadda_tree_6(2)(11);
	dadda_tree_5(3)(11) <= dadda_tree_6(3)(11);
	dadda_tree_5(4)(11) <= dadda_tree_6(4)(11);
	dadda_tree_5(5)(11) <= dadda_tree_6(5)(11);
	dadda_tree_5(0)(12) <= dadda_tree_6(0)(12);
	dadda_tree_5(1)(12) <= dadda_tree_6(1)(12);
	dadda_tree_5(2)(12) <= dadda_tree_6(2)(12);
	dadda_tree_5(3)(12) <= dadda_tree_6(3)(12);
	dadda_tree_5(4)(12) <= dadda_tree_6(4)(12);
	dadda_tree_5(5)(12) <= dadda_tree_6(5)(12);
	dadda_tree_5(6)(12) <= dadda_tree_6(6)(12);
	dadda_tree_5(7)(12) <= dadda_tree_6(7)(12);
	dadda_tree_5(0)(13) <= dadda_tree_6(0)(13);
	dadda_tree_5(1)(13) <= dadda_tree_6(1)(13);
	dadda_tree_5(2)(13) <= dadda_tree_6(2)(13);
	dadda_tree_5(3)(13) <= dadda_tree_6(3)(13);
	dadda_tree_5(4)(13) <= dadda_tree_6(4)(13);
	dadda_tree_5(5)(13) <= dadda_tree_6(5)(13);
	dadda_tree_5(6)(13) <= dadda_tree_6(6)(13);
	dadda_tree_5(0)(14) <= dadda_tree_6(0)(14);
	dadda_tree_5(1)(14) <= dadda_tree_6(1)(14);
	dadda_tree_5(2)(14) <= dadda_tree_6(2)(14);
	dadda_tree_5(3)(14) <= dadda_tree_6(3)(14);
	dadda_tree_5(4)(14) <= dadda_tree_6(4)(14);
	dadda_tree_5(5)(14) <= dadda_tree_6(5)(14);
	dadda_tree_5(6)(14) <= dadda_tree_6(6)(14);
	dadda_tree_5(7)(14) <= dadda_tree_6(7)(14);
	dadda_tree_5(8)(14) <= dadda_tree_6(8)(14);
	dadda_tree_5(0)(15) <= dadda_tree_6(0)(15);
	dadda_tree_5(1)(15) <= dadda_tree_6(1)(15);
	dadda_tree_5(2)(15) <= dadda_tree_6(2)(15);
	dadda_tree_5(3)(15) <= dadda_tree_6(3)(15);
	dadda_tree_5(4)(15) <= dadda_tree_6(4)(15);
	dadda_tree_5(5)(15) <= dadda_tree_6(5)(15);
	dadda_tree_5(6)(15) <= dadda_tree_6(6)(15);
	dadda_tree_5(7)(15) <= dadda_tree_6(7)(15);
	dadda_tree_5(0)(16) <= dadda_tree_6(0)(16);
	dadda_tree_5(1)(16) <= dadda_tree_6(1)(16);
	dadda_tree_5(2)(16) <= dadda_tree_6(2)(16);
	dadda_tree_5(3)(16) <= dadda_tree_6(3)(16);
	dadda_tree_5(4)(16) <= dadda_tree_6(4)(16);
	dadda_tree_5(5)(16) <= dadda_tree_6(5)(16);
	dadda_tree_5(6)(16) <= dadda_tree_6(6)(16);
	dadda_tree_5(7)(16) <= dadda_tree_6(7)(16);
	dadda_tree_5(8)(16) <= dadda_tree_6(8)(16);
	dadda_tree_5(9)(16) <= dadda_tree_6(9)(16);
	dadda_tree_5(0)(17) <= dadda_tree_6(0)(17);
	dadda_tree_5(1)(17) <= dadda_tree_6(1)(17);
	dadda_tree_5(2)(17) <= dadda_tree_6(2)(17);
	dadda_tree_5(3)(17) <= dadda_tree_6(3)(17);
	dadda_tree_5(4)(17) <= dadda_tree_6(4)(17);
	dadda_tree_5(5)(17) <= dadda_tree_6(5)(17);
	dadda_tree_5(6)(17) <= dadda_tree_6(6)(17);
	dadda_tree_5(7)(17) <= dadda_tree_6(7)(17);
	dadda_tree_5(8)(17) <= dadda_tree_6(8)(17);
	dadda_tree_5(0)(18) <= dadda_tree_6(0)(18);
	dadda_tree_5(1)(18) <= dadda_tree_6(1)(18);
	dadda_tree_5(2)(18) <= dadda_tree_6(2)(18);
	dadda_tree_5(3)(18) <= dadda_tree_6(3)(18);
	dadda_tree_5(4)(18) <= dadda_tree_6(4)(18);
	dadda_tree_5(5)(18) <= dadda_tree_6(5)(18);
	dadda_tree_5(6)(18) <= dadda_tree_6(6)(18);
	dadda_tree_5(7)(18) <= dadda_tree_6(7)(18);
	dadda_tree_5(8)(18) <= dadda_tree_6(8)(18);
	dadda_tree_5(9)(18) <= dadda_tree_6(9)(18);
	dadda_tree_5(10)(18) <= dadda_tree_6(10)(18);
	dadda_tree_5(0)(19) <= dadda_tree_6(0)(19);
	dadda_tree_5(1)(19) <= dadda_tree_6(1)(19);
	dadda_tree_5(2)(19) <= dadda_tree_6(2)(19);
	dadda_tree_5(3)(19) <= dadda_tree_6(3)(19);
	dadda_tree_5(4)(19) <= dadda_tree_6(4)(19);
	dadda_tree_5(5)(19) <= dadda_tree_6(5)(19);
	dadda_tree_5(6)(19) <= dadda_tree_6(6)(19);
	dadda_tree_5(7)(19) <= dadda_tree_6(7)(19);
	dadda_tree_5(8)(19) <= dadda_tree_6(8)(19);
	dadda_tree_5(9)(19) <= dadda_tree_6(9)(19);
	dadda_tree_5(0)(20) <= dadda_tree_6(0)(20);
	dadda_tree_5(1)(20) <= dadda_tree_6(1)(20);
	dadda_tree_5(2)(20) <= dadda_tree_6(2)(20);
	dadda_tree_5(3)(20) <= dadda_tree_6(3)(20);
	dadda_tree_5(4)(20) <= dadda_tree_6(4)(20);
	dadda_tree_5(5)(20) <= dadda_tree_6(5)(20);
	dadda_tree_5(6)(20) <= dadda_tree_6(6)(20);
	dadda_tree_5(7)(20) <= dadda_tree_6(7)(20);
	dadda_tree_5(8)(20) <= dadda_tree_6(8)(20);
	dadda_tree_5(9)(20) <= dadda_tree_6(9)(20);
	dadda_tree_5(10)(20) <= dadda_tree_6(10)(20);
	dadda_tree_5(11)(20) <= dadda_tree_6(11)(20);
	dadda_tree_5(0)(21) <= dadda_tree_6(0)(21);
	dadda_tree_5(1)(21) <= dadda_tree_6(1)(21);
	dadda_tree_5(2)(21) <= dadda_tree_6(2)(21);
	dadda_tree_5(3)(21) <= dadda_tree_6(3)(21);
	dadda_tree_5(4)(21) <= dadda_tree_6(4)(21);
	dadda_tree_5(5)(21) <= dadda_tree_6(5)(21);
	dadda_tree_5(6)(21) <= dadda_tree_6(6)(21);
	dadda_tree_5(7)(21) <= dadda_tree_6(7)(21);
	dadda_tree_5(8)(21) <= dadda_tree_6(8)(21);
	dadda_tree_5(9)(21) <= dadda_tree_6(9)(21);
	dadda_tree_5(10)(21) <= dadda_tree_6(10)(21);
	dadda_tree_5(0)(22) <= dadda_tree_6(0)(22);
	dadda_tree_5(1)(22) <= dadda_tree_6(1)(22);
	dadda_tree_5(2)(22) <= dadda_tree_6(2)(22);
	dadda_tree_5(3)(22) <= dadda_tree_6(3)(22);
	dadda_tree_5(4)(22) <= dadda_tree_6(4)(22);
	dadda_tree_5(5)(22) <= dadda_tree_6(5)(22);
	dadda_tree_5(6)(22) <= dadda_tree_6(6)(22);
	dadda_tree_5(7)(22) <= dadda_tree_6(7)(22);
	dadda_tree_5(8)(22) <= dadda_tree_6(8)(22);
	dadda_tree_5(9)(22) <= dadda_tree_6(9)(22);
	dadda_tree_5(10)(22) <= dadda_tree_6(10)(22);
	dadda_tree_5(11)(22) <= dadda_tree_6(11)(22);
	dadda_tree_5(12)(22) <= dadda_tree_6(12)(22);
	dadda_tree_5(0)(23) <= dadda_tree_6(0)(23);
	dadda_tree_5(1)(23) <= dadda_tree_6(1)(23);
	dadda_tree_5(2)(23) <= dadda_tree_6(2)(23);
	dadda_tree_5(3)(23) <= dadda_tree_6(3)(23);
	dadda_tree_5(4)(23) <= dadda_tree_6(4)(23);
	dadda_tree_5(5)(23) <= dadda_tree_6(5)(23);
	dadda_tree_5(6)(23) <= dadda_tree_6(6)(23);
	dadda_tree_5(7)(23) <= dadda_tree_6(7)(23);
	dadda_tree_5(8)(23) <= dadda_tree_6(8)(23);
	dadda_tree_5(9)(23) <= dadda_tree_6(9)(23);
	dadda_tree_5(10)(23) <= dadda_tree_6(10)(23);
	dadda_tree_5(11)(23) <= dadda_tree_6(11)(23);

	ha_6_0_24: ha
		port map(
			a => dadda_tree_6(0)(24),
			b => dadda_tree_6(1)(24),
			s => dadda_tree_5(0)(24),
			co => dadda_tree_5(0)(25)
	);

	dadda_tree_5(1)(24) <= dadda_tree_6(2)(24);
	dadda_tree_5(2)(24) <= dadda_tree_6(3)(24);
	dadda_tree_5(3)(24) <= dadda_tree_6(4)(24);
	dadda_tree_5(4)(24) <= dadda_tree_6(5)(24);
	dadda_tree_5(5)(24) <= dadda_tree_6(6)(24);
	dadda_tree_5(6)(24) <= dadda_tree_6(7)(24);
	dadda_tree_5(7)(24) <= dadda_tree_6(8)(24);
	dadda_tree_5(8)(24) <= dadda_tree_6(9)(24);
	dadda_tree_5(9)(24) <= dadda_tree_6(10)(24);
	dadda_tree_5(10)(24) <= dadda_tree_6(11)(24);
	dadda_tree_5(11)(24) <= dadda_tree_6(12)(24);
	dadda_tree_5(12)(24) <= dadda_tree_6(13)(24);

	ha_6_0_25: ha
		port map(
			a => dadda_tree_6(0)(25),
			b => dadda_tree_6(1)(25),
			s => dadda_tree_5(1)(25),
			co => dadda_tree_5(0)(26)
	);

	dadda_tree_5(2)(25) <= dadda_tree_6(2)(25);
	dadda_tree_5(3)(25) <= dadda_tree_6(3)(25);
	dadda_tree_5(4)(25) <= dadda_tree_6(4)(25);
	dadda_tree_5(5)(25) <= dadda_tree_6(5)(25);
	dadda_tree_5(6)(25) <= dadda_tree_6(6)(25);
	dadda_tree_5(7)(25) <= dadda_tree_6(7)(25);
	dadda_tree_5(8)(25) <= dadda_tree_6(8)(25);
	dadda_tree_5(9)(25) <= dadda_tree_6(9)(25);
	dadda_tree_5(10)(25) <= dadda_tree_6(10)(25);
	dadda_tree_5(11)(25) <= dadda_tree_6(11)(25);
	dadda_tree_5(12)(25) <= dadda_tree_6(12)(25);

	fa_6_0_26: fa
		port map(
			a => dadda_tree_6(0)(26),
			b => dadda_tree_6(1)(26),
			ci => dadda_tree_6(2)(26),
			s => dadda_tree_5(1)(26),
			co => dadda_tree_5(0)(27)
	);

	ha_6_3_26: ha
		port map(
			a => dadda_tree_6(3)(26),
			b => dadda_tree_6(4)(26),
			s => dadda_tree_5(2)(26),
			co => dadda_tree_5(1)(27)
	);

	dadda_tree_5(3)(26) <= dadda_tree_6(5)(26);
	dadda_tree_5(4)(26) <= dadda_tree_6(6)(26);
	dadda_tree_5(5)(26) <= dadda_tree_6(7)(26);
	dadda_tree_5(6)(26) <= dadda_tree_6(8)(26);
	dadda_tree_5(7)(26) <= dadda_tree_6(9)(26);
	dadda_tree_5(8)(26) <= dadda_tree_6(10)(26);
	dadda_tree_5(9)(26) <= dadda_tree_6(11)(26);
	dadda_tree_5(10)(26) <= dadda_tree_6(12)(26);
	dadda_tree_5(11)(26) <= dadda_tree_6(13)(26);
	dadda_tree_5(12)(26) <= dadda_tree_6(14)(26);

	fa_6_0_27: fa
		port map(
			a => dadda_tree_6(0)(27),
			b => dadda_tree_6(1)(27),
			ci => dadda_tree_6(2)(27),
			s => dadda_tree_5(2)(27),
			co => dadda_tree_5(0)(28)
	);

	ha_6_3_27: ha
		port map(
			a => dadda_tree_6(3)(27),
			b => dadda_tree_6(4)(27),
			s => dadda_tree_5(3)(27),
			co => dadda_tree_5(1)(28)
	);

	dadda_tree_5(4)(27) <= dadda_tree_6(5)(27);
	dadda_tree_5(5)(27) <= dadda_tree_6(6)(27);
	dadda_tree_5(6)(27) <= dadda_tree_6(7)(27);
	dadda_tree_5(7)(27) <= dadda_tree_6(8)(27);
	dadda_tree_5(8)(27) <= dadda_tree_6(9)(27);
	dadda_tree_5(9)(27) <= dadda_tree_6(10)(27);
	dadda_tree_5(10)(27) <= dadda_tree_6(11)(27);
	dadda_tree_5(11)(27) <= dadda_tree_6(12)(27);
	dadda_tree_5(12)(27) <= dadda_tree_6(13)(27);

	fa_6_0_28: fa
		port map(
			a => dadda_tree_6(0)(28),
			b => dadda_tree_6(1)(28),
			ci => dadda_tree_6(2)(28),
			s => dadda_tree_5(2)(28),
			co => dadda_tree_5(0)(29)
	);

	fa_6_3_28: fa
		port map(
			a => dadda_tree_6(3)(28),
			b => dadda_tree_6(4)(28),
			ci => dadda_tree_6(5)(28),
			s => dadda_tree_5(3)(28),
			co => dadda_tree_5(1)(29)
	);

	ha_6_6_28: ha
		port map(
			a => dadda_tree_6(6)(28),
			b => dadda_tree_6(7)(28),
			s => dadda_tree_5(4)(28),
			co => dadda_tree_5(2)(29)
	);

	dadda_tree_5(5)(28) <= dadda_tree_6(8)(28);
	dadda_tree_5(6)(28) <= dadda_tree_6(9)(28);
	dadda_tree_5(7)(28) <= dadda_tree_6(10)(28);
	dadda_tree_5(8)(28) <= dadda_tree_6(11)(28);
	dadda_tree_5(9)(28) <= dadda_tree_6(12)(28);
	dadda_tree_5(10)(28) <= dadda_tree_6(13)(28);
	dadda_tree_5(11)(28) <= dadda_tree_6(14)(28);
	dadda_tree_5(12)(28) <= dadda_tree_6(15)(28);

	fa_6_0_29: fa
		port map(
			a => dadda_tree_6(0)(29),
			b => dadda_tree_6(1)(29),
			ci => dadda_tree_6(2)(29),
			s => dadda_tree_5(3)(29),
			co => dadda_tree_5(0)(30)
	);

	fa_6_3_29: fa
		port map(
			a => dadda_tree_6(3)(29),
			b => dadda_tree_6(4)(29),
			ci => dadda_tree_6(5)(29),
			s => dadda_tree_5(4)(29),
			co => dadda_tree_5(1)(30)
	);

	ha_6_6_29: ha
		port map(
			a => dadda_tree_6(6)(29),
			b => dadda_tree_6(7)(29),
			s => dadda_tree_5(5)(29),
			co => dadda_tree_5(2)(30)
	);

	dadda_tree_5(6)(29) <= dadda_tree_6(8)(29);
	dadda_tree_5(7)(29) <= dadda_tree_6(9)(29);
	dadda_tree_5(8)(29) <= dadda_tree_6(10)(29);
	dadda_tree_5(9)(29) <= dadda_tree_6(11)(29);
	dadda_tree_5(10)(29) <= dadda_tree_6(12)(29);
	dadda_tree_5(11)(29) <= dadda_tree_6(13)(29);
	dadda_tree_5(12)(29) <= dadda_tree_6(14)(29);

	fa_6_0_30: fa
		port map(
			a => dadda_tree_6(0)(30),
			b => dadda_tree_6(1)(30),
			ci => dadda_tree_6(2)(30),
			s => dadda_tree_5(3)(30),
			co => dadda_tree_5(0)(31)
	);

	fa_6_3_30: fa
		port map(
			a => dadda_tree_6(3)(30),
			b => dadda_tree_6(4)(30),
			ci => dadda_tree_6(5)(30),
			s => dadda_tree_5(4)(30),
			co => dadda_tree_5(1)(31)
	);

	fa_6_6_30: fa
		port map(
			a => dadda_tree_6(6)(30),
			b => dadda_tree_6(7)(30),
			ci => dadda_tree_6(8)(30),
			s => dadda_tree_5(5)(30),
			co => dadda_tree_5(2)(31)
	);

	ha_6_9_30: ha
		port map(
			a => dadda_tree_6(9)(30),
			b => dadda_tree_6(10)(30),
			s => dadda_tree_5(6)(30),
			co => dadda_tree_5(3)(31)
	);

	dadda_tree_5(7)(30) <= dadda_tree_6(11)(30);
	dadda_tree_5(8)(30) <= dadda_tree_6(12)(30);
	dadda_tree_5(9)(30) <= dadda_tree_6(13)(30);
	dadda_tree_5(10)(30) <= dadda_tree_6(14)(30);
	dadda_tree_5(11)(30) <= dadda_tree_6(15)(30);
	dadda_tree_5(12)(30) <= dadda_tree_6(16)(30);

	fa_6_0_31: fa
		port map(
			a => dadda_tree_6(0)(31),
			b => dadda_tree_6(1)(31),
			ci => dadda_tree_6(2)(31),
			s => dadda_tree_5(4)(31),
			co => dadda_tree_5(0)(32)
	);

	fa_6_3_31: fa
		port map(
			a => dadda_tree_6(3)(31),
			b => dadda_tree_6(4)(31),
			ci => dadda_tree_6(5)(31),
			s => dadda_tree_5(5)(31),
			co => dadda_tree_5(1)(32)
	);

	fa_6_6_31: fa
		port map(
			a => dadda_tree_6(6)(31),
			b => dadda_tree_6(7)(31),
			ci => dadda_tree_6(8)(31),
			s => dadda_tree_5(6)(31),
			co => dadda_tree_5(2)(32)
	);

	ha_6_9_31: ha
		port map(
			a => dadda_tree_6(9)(31),
			b => dadda_tree_6(10)(31),
			s => dadda_tree_5(7)(31),
			co => dadda_tree_5(3)(32)
	);

	dadda_tree_5(8)(31) <= dadda_tree_6(11)(31);
	dadda_tree_5(9)(31) <= dadda_tree_6(12)(31);
	dadda_tree_5(10)(31) <= dadda_tree_6(13)(31);
	dadda_tree_5(11)(31) <= dadda_tree_6(14)(31);
	dadda_tree_5(12)(31) <= dadda_tree_6(15)(31);

	fa_6_0_32: fa
		port map(
			a => dadda_tree_6(0)(32),
			b => dadda_tree_6(1)(32),
			ci => dadda_tree_6(2)(32),
			s => dadda_tree_5(4)(32),
			co => dadda_tree_5(0)(33)
	);

	fa_6_3_32: fa
		port map(
			a => dadda_tree_6(3)(32),
			b => dadda_tree_6(4)(32),
			ci => dadda_tree_6(5)(32),
			s => dadda_tree_5(5)(32),
			co => dadda_tree_5(1)(33)
	);

	fa_6_6_32: fa
		port map(
			a => dadda_tree_6(6)(32),
			b => dadda_tree_6(7)(32),
			ci => dadda_tree_6(8)(32),
			s => dadda_tree_5(6)(32),
			co => dadda_tree_5(2)(33)
	);

	fa_6_9_32: fa
		port map(
			a => dadda_tree_6(9)(32),
			b => dadda_tree_6(10)(32),
			ci => dadda_tree_6(11)(32),
			s => dadda_tree_5(7)(32),
			co => dadda_tree_5(3)(33)
	);
	dadda_tree_5(8)(32) <= dadda_tree_6(12)(32);
	dadda_tree_5(9)(32) <= dadda_tree_6(13)(32);
	dadda_tree_5(10)(32) <= dadda_tree_6(14)(32);
	dadda_tree_5(11)(32) <= dadda_tree_6(15)(32);
	dadda_tree_5(12)(32) <= dadda_tree_6(16)(32);

	fa_6_0_33: fa
		port map(
			a => dadda_tree_6(0)(33),
			b => dadda_tree_6(1)(33),
			ci => dadda_tree_6(2)(33),
			s => dadda_tree_5(4)(33),
			co => dadda_tree_5(0)(34)
	);

	fa_6_3_33: fa
		port map(
			a => dadda_tree_6(3)(33),
			b => dadda_tree_6(4)(33),
			ci => dadda_tree_6(5)(33),
			s => dadda_tree_5(5)(33),
			co => dadda_tree_5(1)(34)
	);

	fa_6_6_33: fa
		port map(
			a => dadda_tree_6(6)(33),
			b => dadda_tree_6(7)(33),
			ci => dadda_tree_6(8)(33),
			s => dadda_tree_5(6)(33),
			co => dadda_tree_5(2)(34)
	);

	fa_6_9_33: fa
		port map(
			a => dadda_tree_6(9)(33),
			b => dadda_tree_6(10)(33),
			ci => dadda_tree_6(11)(33),
			s => dadda_tree_5(7)(33),
			co => dadda_tree_5(3)(34)
	);
	dadda_tree_5(8)(33) <= dadda_tree_6(12)(33);
	dadda_tree_5(9)(33) <= dadda_tree_6(13)(33);
	dadda_tree_5(10)(33) <= dadda_tree_6(14)(33);
	dadda_tree_5(11)(33) <= dadda_tree_6(15)(33);
	dadda_tree_5(12)(33) <= dadda_tree_6(16)(33);

	fa_6_0_34: fa
		port map(
			a => dadda_tree_6(0)(34),
			b => dadda_tree_6(1)(34),
			ci => dadda_tree_6(2)(34),
			s => dadda_tree_5(4)(34),
			co => dadda_tree_5(0)(35)
	);

	fa_6_3_34: fa
		port map(
			a => dadda_tree_6(3)(34),
			b => dadda_tree_6(4)(34),
			ci => dadda_tree_6(5)(34),
			s => dadda_tree_5(5)(34),
			co => dadda_tree_5(1)(35)
	);

	fa_6_6_34: fa
		port map(
			a => dadda_tree_6(6)(34),
			b => dadda_tree_6(7)(34),
			ci => dadda_tree_6(8)(34),
			s => dadda_tree_5(6)(34),
			co => dadda_tree_5(2)(35)
	);

	fa_6_9_34: fa
		port map(
			a => dadda_tree_6(9)(34),
			b => dadda_tree_6(10)(34),
			ci => dadda_tree_6(11)(34),
			s => dadda_tree_5(7)(34),
			co => dadda_tree_5(3)(35)
	);
	dadda_tree_5(8)(34) <= dadda_tree_6(12)(34);
	dadda_tree_5(9)(34) <= dadda_tree_6(13)(34);
	dadda_tree_5(10)(34) <= dadda_tree_6(14)(34);
	dadda_tree_5(11)(34) <= dadda_tree_6(15)(34);
	dadda_tree_5(12)(34) <= dadda_tree_6(16)(34);

	fa_6_0_35: fa
		port map(
			a => dadda_tree_6(0)(35),
			b => dadda_tree_6(1)(35),
			ci => dadda_tree_6(2)(35),
			s => dadda_tree_5(4)(35),
			co => dadda_tree_5(0)(36)
	);

	fa_6_3_35: fa
		port map(
			a => dadda_tree_6(3)(35),
			b => dadda_tree_6(4)(35),
			ci => dadda_tree_6(5)(35),
			s => dadda_tree_5(5)(35),
			co => dadda_tree_5(1)(36)
	);

	fa_6_6_35: fa
		port map(
			a => dadda_tree_6(6)(35),
			b => dadda_tree_6(7)(35),
			ci => dadda_tree_6(8)(35),
			s => dadda_tree_5(6)(35),
			co => dadda_tree_5(2)(36)
	);

	fa_6_9_35: fa
		port map(
			a => dadda_tree_6(9)(35),
			b => dadda_tree_6(10)(35),
			ci => dadda_tree_6(11)(35),
			s => dadda_tree_5(7)(35),
			co => dadda_tree_5(3)(36)
	);
	dadda_tree_5(8)(35) <= dadda_tree_6(12)(35);
	dadda_tree_5(9)(35) <= dadda_tree_6(13)(35);
	dadda_tree_5(10)(35) <= dadda_tree_6(14)(35);
	dadda_tree_5(11)(35) <= dadda_tree_6(15)(35);
	dadda_tree_5(12)(35) <= dadda_tree_6(16)(35);

	fa_6_1_36: fa
		port map(
			a => dadda_tree_6(1)(36),
			b => dadda_tree_6(2)(36),
			ci => dadda_tree_6(3)(36),
			s => dadda_tree_5(4)(36),
			co => dadda_tree_5(0)(37)
	);

	fa_6_4_36: fa
		port map(
			a => dadda_tree_6(4)(36),
			b => dadda_tree_6(5)(36),
			ci => dadda_tree_6(6)(36),
			s => dadda_tree_5(5)(36),
			co => dadda_tree_5(1)(37)
	);

	fa_6_7_36: fa
		port map(
			a => dadda_tree_6(7)(36),
			b => dadda_tree_6(8)(36),
			ci => dadda_tree_6(9)(36),
			s => dadda_tree_5(6)(36),
			co => dadda_tree_5(2)(37)
	);

	ha_6_10_36: ha
		port map(
			a => dadda_tree_6(10)(36),
			b => dadda_tree_6(11)(36),
			s => dadda_tree_5(7)(36),
			co => dadda_tree_5(3)(37)
	);

	dadda_tree_5(8)(36) <= dadda_tree_6(12)(36);
	dadda_tree_5(9)(36) <= dadda_tree_6(13)(36);
	dadda_tree_5(10)(36) <= dadda_tree_6(14)(36);
	dadda_tree_5(11)(36) <= dadda_tree_6(15)(36);
	dadda_tree_5(12)(36) <= dadda_tree_6(16)(36);

	fa_6_2_37: fa
		port map(
			a => dadda_tree_6(2)(37),
			b => dadda_tree_6(3)(37),
			ci => dadda_tree_6(4)(37),
			s => dadda_tree_5(4)(37),
			co => dadda_tree_5(0)(38)
	);

	fa_6_5_37: fa
		port map(
			a => dadda_tree_6(5)(37),
			b => dadda_tree_6(6)(37),
			ci => dadda_tree_6(7)(37),
			s => dadda_tree_5(5)(37),
			co => dadda_tree_5(1)(38)
	);

	fa_6_8_37: fa
		port map(
			a => dadda_tree_6(8)(37),
			b => dadda_tree_6(9)(37),
			ci => dadda_tree_6(10)(37),
			s => dadda_tree_5(6)(37),
			co => dadda_tree_5(2)(38)
	);
	dadda_tree_5(7)(37) <= dadda_tree_6(11)(37);
	dadda_tree_5(8)(37) <= dadda_tree_6(12)(37);
	dadda_tree_5(9)(37) <= dadda_tree_6(13)(37);
	dadda_tree_5(10)(37) <= dadda_tree_6(14)(37);
	dadda_tree_5(11)(37) <= dadda_tree_6(15)(37);
	dadda_tree_5(12)(37) <= dadda_tree_6(16)(37);

	fa_6_2_38: fa
		port map(
			a => dadda_tree_6(2)(38),
			b => dadda_tree_6(3)(38),
			ci => dadda_tree_6(4)(38),
			s => dadda_tree_5(3)(38),
			co => dadda_tree_5(0)(39)
	);

	fa_6_5_38: fa
		port map(
			a => dadda_tree_6(5)(38),
			b => dadda_tree_6(6)(38),
			ci => dadda_tree_6(7)(38),
			s => dadda_tree_5(4)(38),
			co => dadda_tree_5(1)(39)
	);

	ha_6_8_38: ha
		port map(
			a => dadda_tree_6(8)(38),
			b => dadda_tree_6(9)(38),
			s => dadda_tree_5(5)(38),
			co => dadda_tree_5(2)(39)
	);

	dadda_tree_5(6)(38) <= dadda_tree_6(10)(38);
	dadda_tree_5(7)(38) <= dadda_tree_6(11)(38);
	dadda_tree_5(8)(38) <= dadda_tree_6(12)(38);
	dadda_tree_5(9)(38) <= dadda_tree_6(13)(38);
	dadda_tree_5(10)(38) <= dadda_tree_6(14)(38);
	dadda_tree_5(11)(38) <= dadda_tree_6(15)(38);
	dadda_tree_5(12)(38) <= dadda_tree_6(16)(38);

	fa_6_3_39: fa
		port map(
			a => dadda_tree_6(3)(39),
			b => dadda_tree_6(4)(39),
			ci => dadda_tree_6(5)(39),
			s => dadda_tree_5(3)(39),
			co => dadda_tree_5(0)(40)
	);

	fa_6_6_39: fa
		port map(
			a => dadda_tree_6(6)(39),
			b => dadda_tree_6(7)(39),
			ci => dadda_tree_6(8)(39),
			s => dadda_tree_5(4)(39),
			co => dadda_tree_5(1)(40)
	);
	dadda_tree_5(5)(39) <= dadda_tree_6(9)(39);
	dadda_tree_5(6)(39) <= dadda_tree_6(10)(39);
	dadda_tree_5(7)(39) <= dadda_tree_6(11)(39);
	dadda_tree_5(8)(39) <= dadda_tree_6(12)(39);
	dadda_tree_5(9)(39) <= dadda_tree_6(13)(39);
	dadda_tree_5(10)(39) <= dadda_tree_6(14)(39);
	dadda_tree_5(11)(39) <= dadda_tree_6(15)(39);
	dadda_tree_5(12)(39) <= dadda_tree_6(16)(39);

	fa_6_3_40: fa
		port map(
			a => dadda_tree_6(3)(40),
			b => dadda_tree_6(4)(40),
			ci => dadda_tree_6(5)(40),
			s => dadda_tree_5(2)(40),
			co => dadda_tree_5(0)(41)
	);

	ha_6_6_40: ha
		port map(
			a => dadda_tree_6(6)(40),
			b => dadda_tree_6(7)(40),
			s => dadda_tree_5(3)(40),
			co => dadda_tree_5(1)(41)
	);

	dadda_tree_5(4)(40) <= dadda_tree_6(8)(40);
	dadda_tree_5(5)(40) <= dadda_tree_6(9)(40);
	dadda_tree_5(6)(40) <= dadda_tree_6(10)(40);
	dadda_tree_5(7)(40) <= dadda_tree_6(11)(40);
	dadda_tree_5(8)(40) <= dadda_tree_6(12)(40);
	dadda_tree_5(9)(40) <= dadda_tree_6(13)(40);
	dadda_tree_5(10)(40) <= dadda_tree_6(14)(40);
	dadda_tree_5(11)(40) <= dadda_tree_6(15)(40);
	dadda_tree_5(12)(40) <= dadda_tree_6(16)(40);

	fa_6_4_41: fa
		port map(
			a => dadda_tree_6(4)(41),
			b => dadda_tree_6(5)(41),
			ci => dadda_tree_6(6)(41),
			s => dadda_tree_5(2)(41),
			co => dadda_tree_5(0)(42)
	);
	dadda_tree_5(3)(41) <= dadda_tree_6(7)(41);
	dadda_tree_5(4)(41) <= dadda_tree_6(8)(41);
	dadda_tree_5(5)(41) <= dadda_tree_6(9)(41);
	dadda_tree_5(6)(41) <= dadda_tree_6(10)(41);
	dadda_tree_5(7)(41) <= dadda_tree_6(11)(41);
	dadda_tree_5(8)(41) <= dadda_tree_6(12)(41);
	dadda_tree_5(9)(41) <= dadda_tree_6(13)(41);
	dadda_tree_5(10)(41) <= dadda_tree_6(14)(41);
	dadda_tree_5(11)(41) <= dadda_tree_6(15)(41);
	dadda_tree_5(12)(41) <= dadda_tree_6(16)(41);

	ha_6_4_42: ha
		port map(
			a => dadda_tree_6(4)(42),
			b => dadda_tree_6(5)(42),
			s => dadda_tree_5(1)(42),
			co => dadda_tree_5(0)(43)
	);

	dadda_tree_5(2)(42) <= dadda_tree_6(6)(42);
	dadda_tree_5(3)(42) <= dadda_tree_6(7)(42);
	dadda_tree_5(4)(42) <= dadda_tree_6(8)(42);
	dadda_tree_5(5)(42) <= dadda_tree_6(9)(42);
	dadda_tree_5(6)(42) <= dadda_tree_6(10)(42);
	dadda_tree_5(7)(42) <= dadda_tree_6(11)(42);
	dadda_tree_5(8)(42) <= dadda_tree_6(12)(42);
	dadda_tree_5(9)(42) <= dadda_tree_6(13)(42);
	dadda_tree_5(10)(42) <= dadda_tree_6(14)(42);
	dadda_tree_5(11)(42) <= dadda_tree_6(15)(42);
	dadda_tree_5(12)(42) <= dadda_tree_6(16)(42);
	dadda_tree_5(0)(43) <= dadda_tree_6(5)(43);
	dadda_tree_5(1)(43) <= dadda_tree_6(6)(43);
	dadda_tree_5(2)(43) <= dadda_tree_6(7)(43);
	dadda_tree_5(3)(43) <= dadda_tree_6(8)(43);
	dadda_tree_5(4)(43) <= dadda_tree_6(9)(43);
	dadda_tree_5(5)(43) <= dadda_tree_6(10)(43);
	dadda_tree_5(6)(43) <= dadda_tree_6(11)(43);
	dadda_tree_5(7)(43) <= dadda_tree_6(12)(43);
	dadda_tree_5(8)(43) <= dadda_tree_6(13)(43);
	dadda_tree_5(9)(43) <= dadda_tree_6(14)(43);
	dadda_tree_5(10)(43) <= dadda_tree_6(15)(43);
	dadda_tree_5(11)(43) <= dadda_tree_6(16)(43);
	dadda_tree_5(0)(44) <= dadda_tree_6(5)(44);
	dadda_tree_5(1)(44) <= dadda_tree_6(6)(44);
	dadda_tree_5(2)(44) <= dadda_tree_6(7)(44);
	dadda_tree_5(3)(44) <= dadda_tree_6(8)(44);
	dadda_tree_5(4)(44) <= dadda_tree_6(9)(44);
	dadda_tree_5(5)(44) <= dadda_tree_6(10)(44);
	dadda_tree_5(6)(44) <= dadda_tree_6(11)(44);
	dadda_tree_5(7)(44) <= dadda_tree_6(12)(44);
	dadda_tree_5(8)(44) <= dadda_tree_6(13)(44);
	dadda_tree_5(9)(44) <= dadda_tree_6(14)(44);
	dadda_tree_5(10)(44) <= dadda_tree_6(15)(44);
	dadda_tree_5(11)(44) <= dadda_tree_6(16)(44);
	dadda_tree_5(0)(45) <= dadda_tree_6(6)(45);
	dadda_tree_5(1)(45) <= dadda_tree_6(7)(45);
	dadda_tree_5(2)(45) <= dadda_tree_6(8)(45);
	dadda_tree_5(3)(45) <= dadda_tree_6(9)(45);
	dadda_tree_5(4)(45) <= dadda_tree_6(10)(45);
	dadda_tree_5(5)(45) <= dadda_tree_6(11)(45);
	dadda_tree_5(6)(45) <= dadda_tree_6(12)(45);
	dadda_tree_5(7)(45) <= dadda_tree_6(13)(45);
	dadda_tree_5(8)(45) <= dadda_tree_6(14)(45);
	dadda_tree_5(9)(45) <= dadda_tree_6(15)(45);
	dadda_tree_5(10)(45) <= dadda_tree_6(16)(45);
	dadda_tree_5(0)(46) <= dadda_tree_6(6)(46);
	dadda_tree_5(1)(46) <= dadda_tree_6(7)(46);
	dadda_tree_5(2)(46) <= dadda_tree_6(8)(46);
	dadda_tree_5(3)(46) <= dadda_tree_6(9)(46);
	dadda_tree_5(4)(46) <= dadda_tree_6(10)(46);
	dadda_tree_5(5)(46) <= dadda_tree_6(11)(46);
	dadda_tree_5(6)(46) <= dadda_tree_6(12)(46);
	dadda_tree_5(7)(46) <= dadda_tree_6(13)(46);
	dadda_tree_5(8)(46) <= dadda_tree_6(14)(46);
	dadda_tree_5(9)(46) <= dadda_tree_6(15)(46);
	dadda_tree_5(10)(46) <= dadda_tree_6(16)(46);
	dadda_tree_5(0)(47) <= dadda_tree_6(7)(47);
	dadda_tree_5(1)(47) <= dadda_tree_6(8)(47);
	dadda_tree_5(2)(47) <= dadda_tree_6(9)(47);
	dadda_tree_5(3)(47) <= dadda_tree_6(10)(47);
	dadda_tree_5(4)(47) <= dadda_tree_6(11)(47);
	dadda_tree_5(5)(47) <= dadda_tree_6(12)(47);
	dadda_tree_5(6)(47) <= dadda_tree_6(13)(47);
	dadda_tree_5(7)(47) <= dadda_tree_6(14)(47);
	dadda_tree_5(8)(47) <= dadda_tree_6(15)(47);
	dadda_tree_5(9)(47) <= dadda_tree_6(16)(47);
	dadda_tree_5(0)(48) <= dadda_tree_6(7)(48);
	dadda_tree_5(1)(48) <= dadda_tree_6(8)(48);
	dadda_tree_5(2)(48) <= dadda_tree_6(9)(48);
	dadda_tree_5(3)(48) <= dadda_tree_6(10)(48);
	dadda_tree_5(4)(48) <= dadda_tree_6(11)(48);
	dadda_tree_5(5)(48) <= dadda_tree_6(12)(48);
	dadda_tree_5(6)(48) <= dadda_tree_6(13)(48);
	dadda_tree_5(7)(48) <= dadda_tree_6(14)(48);
	dadda_tree_5(8)(48) <= dadda_tree_6(15)(48);
	dadda_tree_5(9)(48) <= dadda_tree_6(16)(48);
	dadda_tree_5(0)(49) <= dadda_tree_6(8)(49);
	dadda_tree_5(1)(49) <= dadda_tree_6(9)(49);
	dadda_tree_5(2)(49) <= dadda_tree_6(10)(49);
	dadda_tree_5(3)(49) <= dadda_tree_6(11)(49);
	dadda_tree_5(4)(49) <= dadda_tree_6(12)(49);
	dadda_tree_5(5)(49) <= dadda_tree_6(13)(49);
	dadda_tree_5(6)(49) <= dadda_tree_6(14)(49);
	dadda_tree_5(7)(49) <= dadda_tree_6(15)(49);
	dadda_tree_5(8)(49) <= dadda_tree_6(16)(49);
	dadda_tree_5(0)(50) <= dadda_tree_6(8)(50);
	dadda_tree_5(1)(50) <= dadda_tree_6(9)(50);
	dadda_tree_5(2)(50) <= dadda_tree_6(10)(50);
	dadda_tree_5(3)(50) <= dadda_tree_6(11)(50);
	dadda_tree_5(4)(50) <= dadda_tree_6(12)(50);
	dadda_tree_5(5)(50) <= dadda_tree_6(13)(50);
	dadda_tree_5(6)(50) <= dadda_tree_6(14)(50);
	dadda_tree_5(7)(50) <= dadda_tree_6(15)(50);
	dadda_tree_5(8)(50) <= dadda_tree_6(16)(50);
	dadda_tree_5(0)(51) <= dadda_tree_6(9)(51);
	dadda_tree_5(1)(51) <= dadda_tree_6(10)(51);
	dadda_tree_5(2)(51) <= dadda_tree_6(11)(51);
	dadda_tree_5(3)(51) <= dadda_tree_6(12)(51);
	dadda_tree_5(4)(51) <= dadda_tree_6(13)(51);
	dadda_tree_5(5)(51) <= dadda_tree_6(14)(51);
	dadda_tree_5(6)(51) <= dadda_tree_6(15)(51);
	dadda_tree_5(7)(51) <= dadda_tree_6(16)(51);
	dadda_tree_5(0)(52) <= dadda_tree_6(9)(52);
	dadda_tree_5(1)(52) <= dadda_tree_6(10)(52);
	dadda_tree_5(2)(52) <= dadda_tree_6(11)(52);
	dadda_tree_5(3)(52) <= dadda_tree_6(12)(52);
	dadda_tree_5(4)(52) <= dadda_tree_6(13)(52);
	dadda_tree_5(5)(52) <= dadda_tree_6(14)(52);
	dadda_tree_5(6)(52) <= dadda_tree_6(15)(52);
	dadda_tree_5(7)(52) <= dadda_tree_6(16)(52);
	dadda_tree_5(0)(53) <= dadda_tree_6(10)(53);
	dadda_tree_5(1)(53) <= dadda_tree_6(11)(53);
	dadda_tree_5(2)(53) <= dadda_tree_6(12)(53);
	dadda_tree_5(3)(53) <= dadda_tree_6(13)(53);
	dadda_tree_5(4)(53) <= dadda_tree_6(14)(53);
	dadda_tree_5(5)(53) <= dadda_tree_6(15)(53);
	dadda_tree_5(6)(53) <= dadda_tree_6(16)(53);
	dadda_tree_5(0)(54) <= dadda_tree_6(10)(54);
	dadda_tree_5(1)(54) <= dadda_tree_6(11)(54);
	dadda_tree_5(2)(54) <= dadda_tree_6(12)(54);
	dadda_tree_5(3)(54) <= dadda_tree_6(13)(54);
	dadda_tree_5(4)(54) <= dadda_tree_6(14)(54);
	dadda_tree_5(5)(54) <= dadda_tree_6(15)(54);
	dadda_tree_5(6)(54) <= dadda_tree_6(16)(54);
	dadda_tree_5(0)(55) <= dadda_tree_6(11)(55);
	dadda_tree_5(1)(55) <= dadda_tree_6(12)(55);
	dadda_tree_5(2)(55) <= dadda_tree_6(13)(55);
	dadda_tree_5(3)(55) <= dadda_tree_6(14)(55);
	dadda_tree_5(4)(55) <= dadda_tree_6(15)(55);
	dadda_tree_5(5)(55) <= dadda_tree_6(16)(55);
	dadda_tree_5(0)(56) <= dadda_tree_6(11)(56);
	dadda_tree_5(1)(56) <= dadda_tree_6(12)(56);
	dadda_tree_5(2)(56) <= dadda_tree_6(13)(56);
	dadda_tree_5(3)(56) <= dadda_tree_6(14)(56);
	dadda_tree_5(4)(56) <= dadda_tree_6(15)(56);
	dadda_tree_5(5)(56) <= dadda_tree_6(16)(56);
	dadda_tree_5(0)(57) <= dadda_tree_6(12)(57);
	dadda_tree_5(1)(57) <= dadda_tree_6(13)(57);
	dadda_tree_5(2)(57) <= dadda_tree_6(14)(57);
	dadda_tree_5(3)(57) <= dadda_tree_6(15)(57);
	dadda_tree_5(4)(57) <= dadda_tree_6(16)(57);
	dadda_tree_5(0)(58) <= dadda_tree_6(12)(58);
	dadda_tree_5(1)(58) <= dadda_tree_6(13)(58);
	dadda_tree_5(2)(58) <= dadda_tree_6(14)(58);
	dadda_tree_5(3)(58) <= dadda_tree_6(15)(58);
	dadda_tree_5(4)(58) <= dadda_tree_6(16)(58);
	dadda_tree_5(0)(59) <= dadda_tree_6(13)(59);
	dadda_tree_5(1)(59) <= dadda_tree_6(14)(59);
	dadda_tree_5(2)(59) <= dadda_tree_6(15)(59);
	dadda_tree_5(3)(59) <= dadda_tree_6(16)(59);
	dadda_tree_5(0)(60) <= dadda_tree_6(13)(60);
	dadda_tree_5(1)(60) <= dadda_tree_6(14)(60);
	dadda_tree_5(2)(60) <= dadda_tree_6(15)(60);
	dadda_tree_5(3)(60) <= dadda_tree_6(16)(60);
	dadda_tree_5(0)(61) <= dadda_tree_6(14)(61);
	dadda_tree_5(1)(61) <= dadda_tree_6(15)(61);
	dadda_tree_5(2)(61) <= dadda_tree_6(16)(61);
	dadda_tree_5(0)(62) <= dadda_tree_6(14)(62);
	dadda_tree_5(1)(62) <= dadda_tree_6(15)(62);
	dadda_tree_5(2)(62) <= dadda_tree_6(16)(62);
	dadda_tree_5(0)(63) <= dadda_tree_6(15)(63);
	dadda_tree_5(1)(63) <= dadda_tree_6(16)(63);
	dadda_tree_4(0)(0) <= dadda_tree_5(0)(0);
	dadda_tree_4(1)(0) <= dadda_tree_5(1)(0);
	dadda_tree_4(0)(1) <= dadda_tree_5(0)(1);
	dadda_tree_4(0)(2) <= dadda_tree_5(0)(2);
	dadda_tree_4(1)(2) <= dadda_tree_5(1)(2);
	dadda_tree_4(2)(2) <= dadda_tree_5(2)(2);
	dadda_tree_4(0)(3) <= dadda_tree_5(0)(3);
	dadda_tree_4(1)(3) <= dadda_tree_5(1)(3);
	dadda_tree_4(0)(4) <= dadda_tree_5(0)(4);
	dadda_tree_4(1)(4) <= dadda_tree_5(1)(4);
	dadda_tree_4(2)(4) <= dadda_tree_5(2)(4);
	dadda_tree_4(3)(4) <= dadda_tree_5(3)(4);
	dadda_tree_4(0)(5) <= dadda_tree_5(0)(5);
	dadda_tree_4(1)(5) <= dadda_tree_5(1)(5);
	dadda_tree_4(2)(5) <= dadda_tree_5(2)(5);
	dadda_tree_4(0)(6) <= dadda_tree_5(0)(6);
	dadda_tree_4(1)(6) <= dadda_tree_5(1)(6);
	dadda_tree_4(2)(6) <= dadda_tree_5(2)(6);
	dadda_tree_4(3)(6) <= dadda_tree_5(3)(6);
	dadda_tree_4(4)(6) <= dadda_tree_5(4)(6);
	dadda_tree_4(0)(7) <= dadda_tree_5(0)(7);
	dadda_tree_4(1)(7) <= dadda_tree_5(1)(7);
	dadda_tree_4(2)(7) <= dadda_tree_5(2)(7);
	dadda_tree_4(3)(7) <= dadda_tree_5(3)(7);
	dadda_tree_4(0)(8) <= dadda_tree_5(0)(8);
	dadda_tree_4(1)(8) <= dadda_tree_5(1)(8);
	dadda_tree_4(2)(8) <= dadda_tree_5(2)(8);
	dadda_tree_4(3)(8) <= dadda_tree_5(3)(8);
	dadda_tree_4(4)(8) <= dadda_tree_5(4)(8);
	dadda_tree_4(5)(8) <= dadda_tree_5(5)(8);
	dadda_tree_4(0)(9) <= dadda_tree_5(0)(9);
	dadda_tree_4(1)(9) <= dadda_tree_5(1)(9);
	dadda_tree_4(2)(9) <= dadda_tree_5(2)(9);
	dadda_tree_4(3)(9) <= dadda_tree_5(3)(9);
	dadda_tree_4(4)(9) <= dadda_tree_5(4)(9);
	dadda_tree_4(0)(10) <= dadda_tree_5(0)(10);
	dadda_tree_4(1)(10) <= dadda_tree_5(1)(10);
	dadda_tree_4(2)(10) <= dadda_tree_5(2)(10);
	dadda_tree_4(3)(10) <= dadda_tree_5(3)(10);
	dadda_tree_4(4)(10) <= dadda_tree_5(4)(10);
	dadda_tree_4(5)(10) <= dadda_tree_5(5)(10);
	dadda_tree_4(6)(10) <= dadda_tree_5(6)(10);
	dadda_tree_4(0)(11) <= dadda_tree_5(0)(11);
	dadda_tree_4(1)(11) <= dadda_tree_5(1)(11);
	dadda_tree_4(2)(11) <= dadda_tree_5(2)(11);
	dadda_tree_4(3)(11) <= dadda_tree_5(3)(11);
	dadda_tree_4(4)(11) <= dadda_tree_5(4)(11);
	dadda_tree_4(5)(11) <= dadda_tree_5(5)(11);
	dadda_tree_4(0)(12) <= dadda_tree_5(0)(12);
	dadda_tree_4(1)(12) <= dadda_tree_5(1)(12);
	dadda_tree_4(2)(12) <= dadda_tree_5(2)(12);
	dadda_tree_4(3)(12) <= dadda_tree_5(3)(12);
	dadda_tree_4(4)(12) <= dadda_tree_5(4)(12);
	dadda_tree_4(5)(12) <= dadda_tree_5(5)(12);
	dadda_tree_4(6)(12) <= dadda_tree_5(6)(12);
	dadda_tree_4(7)(12) <= dadda_tree_5(7)(12);
	dadda_tree_4(0)(13) <= dadda_tree_5(0)(13);
	dadda_tree_4(1)(13) <= dadda_tree_5(1)(13);
	dadda_tree_4(2)(13) <= dadda_tree_5(2)(13);
	dadda_tree_4(3)(13) <= dadda_tree_5(3)(13);
	dadda_tree_4(4)(13) <= dadda_tree_5(4)(13);
	dadda_tree_4(5)(13) <= dadda_tree_5(5)(13);
	dadda_tree_4(6)(13) <= dadda_tree_5(6)(13);
	dadda_tree_4(0)(14) <= dadda_tree_5(0)(14);
	dadda_tree_4(1)(14) <= dadda_tree_5(1)(14);
	dadda_tree_4(2)(14) <= dadda_tree_5(2)(14);
	dadda_tree_4(3)(14) <= dadda_tree_5(3)(14);
	dadda_tree_4(4)(14) <= dadda_tree_5(4)(14);
	dadda_tree_4(5)(14) <= dadda_tree_5(5)(14);
	dadda_tree_4(6)(14) <= dadda_tree_5(6)(14);
	dadda_tree_4(7)(14) <= dadda_tree_5(7)(14);
	dadda_tree_4(8)(14) <= dadda_tree_5(8)(14);
	dadda_tree_4(0)(15) <= dadda_tree_5(0)(15);
	dadda_tree_4(1)(15) <= dadda_tree_5(1)(15);
	dadda_tree_4(2)(15) <= dadda_tree_5(2)(15);
	dadda_tree_4(3)(15) <= dadda_tree_5(3)(15);
	dadda_tree_4(4)(15) <= dadda_tree_5(4)(15);
	dadda_tree_4(5)(15) <= dadda_tree_5(5)(15);
	dadda_tree_4(6)(15) <= dadda_tree_5(6)(15);
	dadda_tree_4(7)(15) <= dadda_tree_5(7)(15);

	ha_5_0_16: ha
		port map(
			a => dadda_tree_5(0)(16),
			b => dadda_tree_5(1)(16),
			s => dadda_tree_4(0)(16),
			co => dadda_tree_4(0)(17)
	);

	dadda_tree_4(1)(16) <= dadda_tree_5(2)(16);
	dadda_tree_4(2)(16) <= dadda_tree_5(3)(16);
	dadda_tree_4(3)(16) <= dadda_tree_5(4)(16);
	dadda_tree_4(4)(16) <= dadda_tree_5(5)(16);
	dadda_tree_4(5)(16) <= dadda_tree_5(6)(16);
	dadda_tree_4(6)(16) <= dadda_tree_5(7)(16);
	dadda_tree_4(7)(16) <= dadda_tree_5(8)(16);
	dadda_tree_4(8)(16) <= dadda_tree_5(9)(16);

	ha_5_0_17: ha
		port map(
			a => dadda_tree_5(0)(17),
			b => dadda_tree_5(1)(17),
			s => dadda_tree_4(1)(17),
			co => dadda_tree_4(0)(18)
	);

	dadda_tree_4(2)(17) <= dadda_tree_5(2)(17);
	dadda_tree_4(3)(17) <= dadda_tree_5(3)(17);
	dadda_tree_4(4)(17) <= dadda_tree_5(4)(17);
	dadda_tree_4(5)(17) <= dadda_tree_5(5)(17);
	dadda_tree_4(6)(17) <= dadda_tree_5(6)(17);
	dadda_tree_4(7)(17) <= dadda_tree_5(7)(17);
	dadda_tree_4(8)(17) <= dadda_tree_5(8)(17);

	fa_5_0_18: fa
		port map(
			a => dadda_tree_5(0)(18),
			b => dadda_tree_5(1)(18),
			ci => dadda_tree_5(2)(18),
			s => dadda_tree_4(1)(18),
			co => dadda_tree_4(0)(19)
	);

	ha_5_3_18: ha
		port map(
			a => dadda_tree_5(3)(18),
			b => dadda_tree_5(4)(18),
			s => dadda_tree_4(2)(18),
			co => dadda_tree_4(1)(19)
	);

	dadda_tree_4(3)(18) <= dadda_tree_5(5)(18);
	dadda_tree_4(4)(18) <= dadda_tree_5(6)(18);
	dadda_tree_4(5)(18) <= dadda_tree_5(7)(18);
	dadda_tree_4(6)(18) <= dadda_tree_5(8)(18);
	dadda_tree_4(7)(18) <= dadda_tree_5(9)(18);
	dadda_tree_4(8)(18) <= dadda_tree_5(10)(18);

	fa_5_0_19: fa
		port map(
			a => dadda_tree_5(0)(19),
			b => dadda_tree_5(1)(19),
			ci => dadda_tree_5(2)(19),
			s => dadda_tree_4(2)(19),
			co => dadda_tree_4(0)(20)
	);

	ha_5_3_19: ha
		port map(
			a => dadda_tree_5(3)(19),
			b => dadda_tree_5(4)(19),
			s => dadda_tree_4(3)(19),
			co => dadda_tree_4(1)(20)
	);

	dadda_tree_4(4)(19) <= dadda_tree_5(5)(19);
	dadda_tree_4(5)(19) <= dadda_tree_5(6)(19);
	dadda_tree_4(6)(19) <= dadda_tree_5(7)(19);
	dadda_tree_4(7)(19) <= dadda_tree_5(8)(19);
	dadda_tree_4(8)(19) <= dadda_tree_5(9)(19);

	fa_5_0_20: fa
		port map(
			a => dadda_tree_5(0)(20),
			b => dadda_tree_5(1)(20),
			ci => dadda_tree_5(2)(20),
			s => dadda_tree_4(2)(20),
			co => dadda_tree_4(0)(21)
	);

	fa_5_3_20: fa
		port map(
			a => dadda_tree_5(3)(20),
			b => dadda_tree_5(4)(20),
			ci => dadda_tree_5(5)(20),
			s => dadda_tree_4(3)(20),
			co => dadda_tree_4(1)(21)
	);

	ha_5_6_20: ha
		port map(
			a => dadda_tree_5(6)(20),
			b => dadda_tree_5(7)(20),
			s => dadda_tree_4(4)(20),
			co => dadda_tree_4(2)(21)
	);

	dadda_tree_4(5)(20) <= dadda_tree_5(8)(20);
	dadda_tree_4(6)(20) <= dadda_tree_5(9)(20);
	dadda_tree_4(7)(20) <= dadda_tree_5(10)(20);
	dadda_tree_4(8)(20) <= dadda_tree_5(11)(20);

	fa_5_0_21: fa
		port map(
			a => dadda_tree_5(0)(21),
			b => dadda_tree_5(1)(21),
			ci => dadda_tree_5(2)(21),
			s => dadda_tree_4(3)(21),
			co => dadda_tree_4(0)(22)
	);

	fa_5_3_21: fa
		port map(
			a => dadda_tree_5(3)(21),
			b => dadda_tree_5(4)(21),
			ci => dadda_tree_5(5)(21),
			s => dadda_tree_4(4)(21),
			co => dadda_tree_4(1)(22)
	);

	ha_5_6_21: ha
		port map(
			a => dadda_tree_5(6)(21),
			b => dadda_tree_5(7)(21),
			s => dadda_tree_4(5)(21),
			co => dadda_tree_4(2)(22)
	);

	dadda_tree_4(6)(21) <= dadda_tree_5(8)(21);
	dadda_tree_4(7)(21) <= dadda_tree_5(9)(21);
	dadda_tree_4(8)(21) <= dadda_tree_5(10)(21);

	fa_5_0_22: fa
		port map(
			a => dadda_tree_5(0)(22),
			b => dadda_tree_5(1)(22),
			ci => dadda_tree_5(2)(22),
			s => dadda_tree_4(3)(22),
			co => dadda_tree_4(0)(23)
	);

	fa_5_3_22: fa
		port map(
			a => dadda_tree_5(3)(22),
			b => dadda_tree_5(4)(22),
			ci => dadda_tree_5(5)(22),
			s => dadda_tree_4(4)(22),
			co => dadda_tree_4(1)(23)
	);

	fa_5_6_22: fa
		port map(
			a => dadda_tree_5(6)(22),
			b => dadda_tree_5(7)(22),
			ci => dadda_tree_5(8)(22),
			s => dadda_tree_4(5)(22),
			co => dadda_tree_4(2)(23)
	);

	ha_5_9_22: ha
		port map(
			a => dadda_tree_5(9)(22),
			b => dadda_tree_5(10)(22),
			s => dadda_tree_4(6)(22),
			co => dadda_tree_4(3)(23)
	);

	dadda_tree_4(7)(22) <= dadda_tree_5(11)(22);
	dadda_tree_4(8)(22) <= dadda_tree_5(12)(22);

	fa_5_0_23: fa
		port map(
			a => dadda_tree_5(0)(23),
			b => dadda_tree_5(1)(23),
			ci => dadda_tree_5(2)(23),
			s => dadda_tree_4(4)(23),
			co => dadda_tree_4(0)(24)
	);

	fa_5_3_23: fa
		port map(
			a => dadda_tree_5(3)(23),
			b => dadda_tree_5(4)(23),
			ci => dadda_tree_5(5)(23),
			s => dadda_tree_4(5)(23),
			co => dadda_tree_4(1)(24)
	);

	fa_5_6_23: fa
		port map(
			a => dadda_tree_5(6)(23),
			b => dadda_tree_5(7)(23),
			ci => dadda_tree_5(8)(23),
			s => dadda_tree_4(6)(23),
			co => dadda_tree_4(2)(24)
	);

	ha_5_9_23: ha
		port map(
			a => dadda_tree_5(9)(23),
			b => dadda_tree_5(10)(23),
			s => dadda_tree_4(7)(23),
			co => dadda_tree_4(3)(24)
	);

	dadda_tree_4(8)(23) <= dadda_tree_5(11)(23);
	dadda_tree_4(0)(24) <= dadda_tree_5(0)(24);
	dadda_tree_4(0)(25) <= dadda_tree_5(0)(25);
	dadda_tree_4(1)(25) <= dadda_tree_5(1)(25);
	dadda_tree_4(0)(26) <= dadda_tree_5(0)(26);
	dadda_tree_4(1)(26) <= dadda_tree_5(1)(26);
	dadda_tree_4(2)(26) <= dadda_tree_5(2)(26);
	dadda_tree_4(0)(27) <= dadda_tree_5(0)(27);
	dadda_tree_4(1)(27) <= dadda_tree_5(1)(27);
	dadda_tree_4(2)(27) <= dadda_tree_5(2)(27);
	dadda_tree_4(3)(27) <= dadda_tree_5(3)(27);
	dadda_tree_4(0)(28) <= dadda_tree_5(0)(28);
	dadda_tree_4(1)(28) <= dadda_tree_5(1)(28);
	dadda_tree_4(2)(28) <= dadda_tree_5(2)(28);
	dadda_tree_4(3)(28) <= dadda_tree_5(3)(28);
	dadda_tree_4(4)(28) <= dadda_tree_5(4)(28);
	dadda_tree_4(0)(29) <= dadda_tree_5(0)(29);
	dadda_tree_4(1)(29) <= dadda_tree_5(1)(29);
	dadda_tree_4(2)(29) <= dadda_tree_5(2)(29);
	dadda_tree_4(3)(29) <= dadda_tree_5(3)(29);
	dadda_tree_4(4)(29) <= dadda_tree_5(4)(29);
	dadda_tree_4(5)(29) <= dadda_tree_5(5)(29);
	dadda_tree_4(0)(30) <= dadda_tree_5(0)(30);
	dadda_tree_4(1)(30) <= dadda_tree_5(1)(30);
	dadda_tree_4(2)(30) <= dadda_tree_5(2)(30);
	dadda_tree_4(3)(30) <= dadda_tree_5(3)(30);
	dadda_tree_4(4)(30) <= dadda_tree_5(4)(30);
	dadda_tree_4(5)(30) <= dadda_tree_5(5)(30);
	dadda_tree_4(6)(30) <= dadda_tree_5(6)(30);
	dadda_tree_4(0)(31) <= dadda_tree_5(0)(31);
	dadda_tree_4(1)(31) <= dadda_tree_5(1)(31);
	dadda_tree_4(2)(31) <= dadda_tree_5(2)(31);
	dadda_tree_4(3)(31) <= dadda_tree_5(3)(31);
	dadda_tree_4(4)(31) <= dadda_tree_5(4)(31);
	dadda_tree_4(5)(31) <= dadda_tree_5(5)(31);
	dadda_tree_4(6)(31) <= dadda_tree_5(6)(31);
	dadda_tree_4(7)(31) <= dadda_tree_5(7)(31);
	dadda_tree_4(0)(32) <= dadda_tree_5(0)(32);
	dadda_tree_4(1)(32) <= dadda_tree_5(1)(32);
	dadda_tree_4(2)(32) <= dadda_tree_5(2)(32);
	dadda_tree_4(3)(32) <= dadda_tree_5(3)(32);
	dadda_tree_4(4)(32) <= dadda_tree_5(4)(32);
	dadda_tree_4(5)(32) <= dadda_tree_5(5)(32);
	dadda_tree_4(6)(32) <= dadda_tree_5(6)(32);
	dadda_tree_4(7)(32) <= dadda_tree_5(7)(32);
	dadda_tree_4(0)(33) <= dadda_tree_5(0)(33);
	dadda_tree_4(1)(33) <= dadda_tree_5(1)(33);
	dadda_tree_4(2)(33) <= dadda_tree_5(2)(33);
	dadda_tree_4(3)(33) <= dadda_tree_5(3)(33);
	dadda_tree_4(4)(33) <= dadda_tree_5(4)(33);
	dadda_tree_4(5)(33) <= dadda_tree_5(5)(33);
	dadda_tree_4(6)(33) <= dadda_tree_5(6)(33);
	dadda_tree_4(7)(33) <= dadda_tree_5(7)(33);
	dadda_tree_4(0)(34) <= dadda_tree_5(0)(34);
	dadda_tree_4(1)(34) <= dadda_tree_5(1)(34);
	dadda_tree_4(2)(34) <= dadda_tree_5(2)(34);
	dadda_tree_4(3)(34) <= dadda_tree_5(3)(34);
	dadda_tree_4(4)(34) <= dadda_tree_5(4)(34);
	dadda_tree_4(5)(34) <= dadda_tree_5(5)(34);
	dadda_tree_4(6)(34) <= dadda_tree_5(6)(34);
	dadda_tree_4(7)(34) <= dadda_tree_5(7)(34);
	dadda_tree_4(0)(35) <= dadda_tree_5(0)(35);
	dadda_tree_4(1)(35) <= dadda_tree_5(1)(35);
	dadda_tree_4(2)(35) <= dadda_tree_5(2)(35);
	dadda_tree_4(3)(35) <= dadda_tree_5(3)(35);
	dadda_tree_4(4)(35) <= dadda_tree_5(4)(35);
	dadda_tree_4(5)(35) <= dadda_tree_5(5)(35);
	dadda_tree_4(6)(35) <= dadda_tree_5(6)(35);
	dadda_tree_4(7)(35) <= dadda_tree_5(7)(35);
	dadda_tree_4(0)(36) <= dadda_tree_5(0)(36);
	dadda_tree_4(1)(36) <= dadda_tree_5(1)(36);
	dadda_tree_4(2)(36) <= dadda_tree_5(2)(36);
	dadda_tree_4(3)(36) <= dadda_tree_5(3)(36);
	dadda_tree_4(4)(36) <= dadda_tree_5(4)(36);
	dadda_tree_4(5)(36) <= dadda_tree_5(5)(36);
	dadda_tree_4(6)(36) <= dadda_tree_5(6)(36);
	dadda_tree_4(7)(36) <= dadda_tree_5(7)(36);
	dadda_tree_4(0)(37) <= dadda_tree_5(0)(37);
	dadda_tree_4(1)(37) <= dadda_tree_5(1)(37);
	dadda_tree_4(2)(37) <= dadda_tree_5(2)(37);
	dadda_tree_4(3)(37) <= dadda_tree_5(3)(37);
	dadda_tree_4(4)(37) <= dadda_tree_5(4)(37);
	dadda_tree_4(5)(37) <= dadda_tree_5(5)(37);
	dadda_tree_4(6)(37) <= dadda_tree_5(6)(37);
	dadda_tree_4(0)(38) <= dadda_tree_5(0)(38);
	dadda_tree_4(1)(38) <= dadda_tree_5(1)(38);
	dadda_tree_4(2)(38) <= dadda_tree_5(2)(38);
	dadda_tree_4(3)(38) <= dadda_tree_5(3)(38);
	dadda_tree_4(4)(38) <= dadda_tree_5(4)(38);
	dadda_tree_4(5)(38) <= dadda_tree_5(5)(38);
	dadda_tree_4(0)(39) <= dadda_tree_5(0)(39);
	dadda_tree_4(1)(39) <= dadda_tree_5(1)(39);
	dadda_tree_4(2)(39) <= dadda_tree_5(2)(39);
	dadda_tree_4(3)(39) <= dadda_tree_5(3)(39);
	dadda_tree_4(4)(39) <= dadda_tree_5(4)(39);
	dadda_tree_4(0)(40) <= dadda_tree_5(0)(40);
	dadda_tree_4(1)(40) <= dadda_tree_5(1)(40);
	dadda_tree_4(2)(40) <= dadda_tree_5(2)(40);
	dadda_tree_4(3)(40) <= dadda_tree_5(3)(40);
	dadda_tree_4(0)(41) <= dadda_tree_5(0)(41);
	dadda_tree_4(1)(41) <= dadda_tree_5(1)(41);
	dadda_tree_4(2)(41) <= dadda_tree_5(2)(41);
	dadda_tree_4(0)(42) <= dadda_tree_5(0)(42);
	dadda_tree_4(1)(42) <= dadda_tree_5(1)(42);

	fa_5_0_43: fa
		port map(
			a => dadda_tree_5(0)(43),
			b => dadda_tree_5(1)(43),
			ci => dadda_tree_5(2)(43),
			s => dadda_tree_4(0)(43),
			co => dadda_tree_4(0)(44)
	);

	ha_5_3_43: ha
		port map(
			a => dadda_tree_5(3)(43),
			b => dadda_tree_5(4)(43),
			s => dadda_tree_4(1)(43),
			co => dadda_tree_4(1)(44)
	);

	dadda_tree_4(2)(43) <= dadda_tree_5(5)(43);
	dadda_tree_4(3)(43) <= dadda_tree_5(6)(43);
	dadda_tree_4(4)(43) <= dadda_tree_5(7)(43);
	dadda_tree_4(5)(43) <= dadda_tree_5(8)(43);
	dadda_tree_4(6)(43) <= dadda_tree_5(9)(43);
	dadda_tree_4(7)(43) <= dadda_tree_5(10)(43);
	dadda_tree_4(8)(43) <= dadda_tree_5(11)(43);

	fa_5_0_44: fa
		port map(
			a => dadda_tree_5(0)(44),
			b => dadda_tree_5(1)(44),
			ci => dadda_tree_5(2)(44),
			s => dadda_tree_4(2)(44),
			co => dadda_tree_4(0)(45)
	);

	fa_5_3_44: fa
		port map(
			a => dadda_tree_5(3)(44),
			b => dadda_tree_5(4)(44),
			ci => dadda_tree_5(5)(44),
			s => dadda_tree_4(3)(44),
			co => dadda_tree_4(1)(45)
	);

	ha_5_6_44: ha
		port map(
			a => dadda_tree_5(6)(44),
			b => dadda_tree_5(7)(44),
			s => dadda_tree_4(4)(44),
			co => dadda_tree_4(2)(45)
	);

	dadda_tree_4(5)(44) <= dadda_tree_5(8)(44);
	dadda_tree_4(6)(44) <= dadda_tree_5(9)(44);
	dadda_tree_4(7)(44) <= dadda_tree_5(10)(44);
	dadda_tree_4(8)(44) <= dadda_tree_5(11)(44);

	fa_5_0_45: fa
		port map(
			a => dadda_tree_5(0)(45),
			b => dadda_tree_5(1)(45),
			ci => dadda_tree_5(2)(45),
			s => dadda_tree_4(3)(45),
			co => dadda_tree_4(0)(46)
	);

	fa_5_3_45: fa
		port map(
			a => dadda_tree_5(3)(45),
			b => dadda_tree_5(4)(45),
			ci => dadda_tree_5(5)(45),
			s => dadda_tree_4(4)(45),
			co => dadda_tree_4(1)(46)
	);

	ha_5_6_45: ha
		port map(
			a => dadda_tree_5(6)(45),
			b => dadda_tree_5(7)(45),
			s => dadda_tree_4(5)(45),
			co => dadda_tree_4(2)(46)
	);

	dadda_tree_4(6)(45) <= dadda_tree_5(8)(45);
	dadda_tree_4(7)(45) <= dadda_tree_5(9)(45);
	dadda_tree_4(8)(45) <= dadda_tree_5(10)(45);

	fa_5_0_46: fa
		port map(
			a => dadda_tree_5(0)(46),
			b => dadda_tree_5(1)(46),
			ci => dadda_tree_5(2)(46),
			s => dadda_tree_4(3)(46),
			co => dadda_tree_4(0)(47)
	);

	fa_5_3_46: fa
		port map(
			a => dadda_tree_5(3)(46),
			b => dadda_tree_5(4)(46),
			ci => dadda_tree_5(5)(46),
			s => dadda_tree_4(4)(46),
			co => dadda_tree_4(1)(47)
	);

	ha_5_6_46: ha
		port map(
			a => dadda_tree_5(6)(46),
			b => dadda_tree_5(7)(46),
			s => dadda_tree_4(5)(46),
			co => dadda_tree_4(2)(47)
	);

	dadda_tree_4(6)(46) <= dadda_tree_5(8)(46);
	dadda_tree_4(7)(46) <= dadda_tree_5(9)(46);
	dadda_tree_4(8)(46) <= dadda_tree_5(10)(46);

	fa_5_0_47: fa
		port map(
			a => dadda_tree_5(0)(47),
			b => dadda_tree_5(1)(47),
			ci => dadda_tree_5(2)(47),
			s => dadda_tree_4(3)(47),
			co => dadda_tree_4(0)(48)
	);

	fa_5_3_47: fa
		port map(
			a => dadda_tree_5(3)(47),
			b => dadda_tree_5(4)(47),
			ci => dadda_tree_5(5)(47),
			s => dadda_tree_4(4)(47),
			co => dadda_tree_4(1)(48)
	);
	dadda_tree_4(5)(47) <= dadda_tree_5(6)(47);
	dadda_tree_4(6)(47) <= dadda_tree_5(7)(47);
	dadda_tree_4(7)(47) <= dadda_tree_5(8)(47);
	dadda_tree_4(8)(47) <= dadda_tree_5(9)(47);

	fa_5_0_48: fa
		port map(
			a => dadda_tree_5(0)(48),
			b => dadda_tree_5(1)(48),
			ci => dadda_tree_5(2)(48),
			s => dadda_tree_4(2)(48),
			co => dadda_tree_4(0)(49)
	);

	ha_5_3_48: ha
		port map(
			a => dadda_tree_5(3)(48),
			b => dadda_tree_5(4)(48),
			s => dadda_tree_4(3)(48),
			co => dadda_tree_4(1)(49)
	);

	dadda_tree_4(4)(48) <= dadda_tree_5(5)(48);
	dadda_tree_4(5)(48) <= dadda_tree_5(6)(48);
	dadda_tree_4(6)(48) <= dadda_tree_5(7)(48);
	dadda_tree_4(7)(48) <= dadda_tree_5(8)(48);
	dadda_tree_4(8)(48) <= dadda_tree_5(9)(48);

	fa_5_0_49: fa
		port map(
			a => dadda_tree_5(0)(49),
			b => dadda_tree_5(1)(49),
			ci => dadda_tree_5(2)(49),
			s => dadda_tree_4(2)(49),
			co => dadda_tree_4(0)(50)
	);
	dadda_tree_4(3)(49) <= dadda_tree_5(3)(49);
	dadda_tree_4(4)(49) <= dadda_tree_5(4)(49);
	dadda_tree_4(5)(49) <= dadda_tree_5(5)(49);
	dadda_tree_4(6)(49) <= dadda_tree_5(6)(49);
	dadda_tree_4(7)(49) <= dadda_tree_5(7)(49);
	dadda_tree_4(8)(49) <= dadda_tree_5(8)(49);

	ha_5_0_50: ha
		port map(
			a => dadda_tree_5(0)(50),
			b => dadda_tree_5(1)(50),
			s => dadda_tree_4(1)(50),
			co => dadda_tree_4(0)(51)
	);

	dadda_tree_4(2)(50) <= dadda_tree_5(2)(50);
	dadda_tree_4(3)(50) <= dadda_tree_5(3)(50);
	dadda_tree_4(4)(50) <= dadda_tree_5(4)(50);
	dadda_tree_4(5)(50) <= dadda_tree_5(5)(50);
	dadda_tree_4(6)(50) <= dadda_tree_5(6)(50);
	dadda_tree_4(7)(50) <= dadda_tree_5(7)(50);
	dadda_tree_4(8)(50) <= dadda_tree_5(8)(50);
	dadda_tree_4(0)(51) <= dadda_tree_5(0)(51);
	dadda_tree_4(1)(51) <= dadda_tree_5(1)(51);
	dadda_tree_4(2)(51) <= dadda_tree_5(2)(51);
	dadda_tree_4(3)(51) <= dadda_tree_5(3)(51);
	dadda_tree_4(4)(51) <= dadda_tree_5(4)(51);
	dadda_tree_4(5)(51) <= dadda_tree_5(5)(51);
	dadda_tree_4(6)(51) <= dadda_tree_5(6)(51);
	dadda_tree_4(7)(51) <= dadda_tree_5(7)(51);
	dadda_tree_4(0)(52) <= dadda_tree_5(0)(52);
	dadda_tree_4(1)(52) <= dadda_tree_5(1)(52);
	dadda_tree_4(2)(52) <= dadda_tree_5(2)(52);
	dadda_tree_4(3)(52) <= dadda_tree_5(3)(52);
	dadda_tree_4(4)(52) <= dadda_tree_5(4)(52);
	dadda_tree_4(5)(52) <= dadda_tree_5(5)(52);
	dadda_tree_4(6)(52) <= dadda_tree_5(6)(52);
	dadda_tree_4(7)(52) <= dadda_tree_5(7)(52);
	dadda_tree_4(0)(53) <= dadda_tree_5(0)(53);
	dadda_tree_4(1)(53) <= dadda_tree_5(1)(53);
	dadda_tree_4(2)(53) <= dadda_tree_5(2)(53);
	dadda_tree_4(3)(53) <= dadda_tree_5(3)(53);
	dadda_tree_4(4)(53) <= dadda_tree_5(4)(53);
	dadda_tree_4(5)(53) <= dadda_tree_5(5)(53);
	dadda_tree_4(6)(53) <= dadda_tree_5(6)(53);
	dadda_tree_4(0)(54) <= dadda_tree_5(0)(54);
	dadda_tree_4(1)(54) <= dadda_tree_5(1)(54);
	dadda_tree_4(2)(54) <= dadda_tree_5(2)(54);
	dadda_tree_4(3)(54) <= dadda_tree_5(3)(54);
	dadda_tree_4(4)(54) <= dadda_tree_5(4)(54);
	dadda_tree_4(5)(54) <= dadda_tree_5(5)(54);
	dadda_tree_4(6)(54) <= dadda_tree_5(6)(54);
	dadda_tree_4(0)(55) <= dadda_tree_5(0)(55);
	dadda_tree_4(1)(55) <= dadda_tree_5(1)(55);
	dadda_tree_4(2)(55) <= dadda_tree_5(2)(55);
	dadda_tree_4(3)(55) <= dadda_tree_5(3)(55);
	dadda_tree_4(4)(55) <= dadda_tree_5(4)(55);
	dadda_tree_4(5)(55) <= dadda_tree_5(5)(55);
	dadda_tree_4(0)(56) <= dadda_tree_5(0)(56);
	dadda_tree_4(1)(56) <= dadda_tree_5(1)(56);
	dadda_tree_4(2)(56) <= dadda_tree_5(2)(56);
	dadda_tree_4(3)(56) <= dadda_tree_5(3)(56);
	dadda_tree_4(4)(56) <= dadda_tree_5(4)(56);
	dadda_tree_4(5)(56) <= dadda_tree_5(5)(56);
	dadda_tree_4(0)(57) <= dadda_tree_5(0)(57);
	dadda_tree_4(1)(57) <= dadda_tree_5(1)(57);
	dadda_tree_4(2)(57) <= dadda_tree_5(2)(57);
	dadda_tree_4(3)(57) <= dadda_tree_5(3)(57);
	dadda_tree_4(4)(57) <= dadda_tree_5(4)(57);
	dadda_tree_4(0)(58) <= dadda_tree_5(0)(58);
	dadda_tree_4(1)(58) <= dadda_tree_5(1)(58);
	dadda_tree_4(2)(58) <= dadda_tree_5(2)(58);
	dadda_tree_4(3)(58) <= dadda_tree_5(3)(58);
	dadda_tree_4(4)(58) <= dadda_tree_5(4)(58);
	dadda_tree_4(0)(59) <= dadda_tree_5(0)(59);
	dadda_tree_4(1)(59) <= dadda_tree_5(1)(59);
	dadda_tree_4(2)(59) <= dadda_tree_5(2)(59);
	dadda_tree_4(3)(59) <= dadda_tree_5(3)(59);
	dadda_tree_4(0)(60) <= dadda_tree_5(0)(60);
	dadda_tree_4(1)(60) <= dadda_tree_5(1)(60);
	dadda_tree_4(2)(60) <= dadda_tree_5(2)(60);
	dadda_tree_4(3)(60) <= dadda_tree_5(3)(60);
	dadda_tree_4(0)(61) <= dadda_tree_5(0)(61);
	dadda_tree_4(1)(61) <= dadda_tree_5(1)(61);
	dadda_tree_4(2)(61) <= dadda_tree_5(2)(61);
	dadda_tree_4(0)(62) <= dadda_tree_5(0)(62);
	dadda_tree_4(1)(62) <= dadda_tree_5(1)(62);
	dadda_tree_4(2)(62) <= dadda_tree_5(2)(62);
	dadda_tree_4(0)(63) <= dadda_tree_5(0)(63);
	dadda_tree_4(1)(63) <= dadda_tree_5(1)(63);
	dadda_tree_3(0)(0) <= dadda_tree_4(0)(0);
	dadda_tree_3(1)(0) <= dadda_tree_4(1)(0);
	dadda_tree_3(0)(1) <= dadda_tree_4(0)(1);
	dadda_tree_3(0)(2) <= dadda_tree_4(0)(2);
	dadda_tree_3(1)(2) <= dadda_tree_4(1)(2);
	dadda_tree_3(2)(2) <= dadda_tree_4(2)(2);
	dadda_tree_3(0)(3) <= dadda_tree_4(0)(3);
	dadda_tree_3(1)(3) <= dadda_tree_4(1)(3);
	dadda_tree_3(0)(4) <= dadda_tree_4(0)(4);
	dadda_tree_3(1)(4) <= dadda_tree_4(1)(4);
	dadda_tree_3(2)(4) <= dadda_tree_4(2)(4);
	dadda_tree_3(3)(4) <= dadda_tree_4(3)(4);
	dadda_tree_3(0)(5) <= dadda_tree_4(0)(5);
	dadda_tree_3(1)(5) <= dadda_tree_4(1)(5);
	dadda_tree_3(2)(5) <= dadda_tree_4(2)(5);
	dadda_tree_3(0)(6) <= dadda_tree_4(0)(6);
	dadda_tree_3(1)(6) <= dadda_tree_4(1)(6);
	dadda_tree_3(2)(6) <= dadda_tree_4(2)(6);
	dadda_tree_3(3)(6) <= dadda_tree_4(3)(6);
	dadda_tree_3(4)(6) <= dadda_tree_4(4)(6);
	dadda_tree_3(0)(7) <= dadda_tree_4(0)(7);
	dadda_tree_3(1)(7) <= dadda_tree_4(1)(7);
	dadda_tree_3(2)(7) <= dadda_tree_4(2)(7);
	dadda_tree_3(3)(7) <= dadda_tree_4(3)(7);
	dadda_tree_3(0)(8) <= dadda_tree_4(0)(8);
	dadda_tree_3(1)(8) <= dadda_tree_4(1)(8);
	dadda_tree_3(2)(8) <= dadda_tree_4(2)(8);
	dadda_tree_3(3)(8) <= dadda_tree_4(3)(8);
	dadda_tree_3(4)(8) <= dadda_tree_4(4)(8);
	dadda_tree_3(5)(8) <= dadda_tree_4(5)(8);
	dadda_tree_3(0)(9) <= dadda_tree_4(0)(9);
	dadda_tree_3(1)(9) <= dadda_tree_4(1)(9);
	dadda_tree_3(2)(9) <= dadda_tree_4(2)(9);
	dadda_tree_3(3)(9) <= dadda_tree_4(3)(9);
	dadda_tree_3(4)(9) <= dadda_tree_4(4)(9);

	ha_4_0_10: ha
		port map(
			a => dadda_tree_4(0)(10),
			b => dadda_tree_4(1)(10),
			s => dadda_tree_3(0)(10),
			co => dadda_tree_3(0)(11)
	);

	dadda_tree_3(1)(10) <= dadda_tree_4(2)(10);
	dadda_tree_3(2)(10) <= dadda_tree_4(3)(10);
	dadda_tree_3(3)(10) <= dadda_tree_4(4)(10);
	dadda_tree_3(4)(10) <= dadda_tree_4(5)(10);
	dadda_tree_3(5)(10) <= dadda_tree_4(6)(10);

	ha_4_0_11: ha
		port map(
			a => dadda_tree_4(0)(11),
			b => dadda_tree_4(1)(11),
			s => dadda_tree_3(1)(11),
			co => dadda_tree_3(0)(12)
	);

	dadda_tree_3(2)(11) <= dadda_tree_4(2)(11);
	dadda_tree_3(3)(11) <= dadda_tree_4(3)(11);
	dadda_tree_3(4)(11) <= dadda_tree_4(4)(11);
	dadda_tree_3(5)(11) <= dadda_tree_4(5)(11);

	fa_4_0_12: fa
		port map(
			a => dadda_tree_4(0)(12),
			b => dadda_tree_4(1)(12),
			ci => dadda_tree_4(2)(12),
			s => dadda_tree_3(1)(12),
			co => dadda_tree_3(0)(13)
	);

	ha_4_3_12: ha
		port map(
			a => dadda_tree_4(3)(12),
			b => dadda_tree_4(4)(12),
			s => dadda_tree_3(2)(12),
			co => dadda_tree_3(1)(13)
	);

	dadda_tree_3(3)(12) <= dadda_tree_4(5)(12);
	dadda_tree_3(4)(12) <= dadda_tree_4(6)(12);
	dadda_tree_3(5)(12) <= dadda_tree_4(7)(12);

	fa_4_0_13: fa
		port map(
			a => dadda_tree_4(0)(13),
			b => dadda_tree_4(1)(13),
			ci => dadda_tree_4(2)(13),
			s => dadda_tree_3(2)(13),
			co => dadda_tree_3(0)(14)
	);

	ha_4_3_13: ha
		port map(
			a => dadda_tree_4(3)(13),
			b => dadda_tree_4(4)(13),
			s => dadda_tree_3(3)(13),
			co => dadda_tree_3(1)(14)
	);

	dadda_tree_3(4)(13) <= dadda_tree_4(5)(13);
	dadda_tree_3(5)(13) <= dadda_tree_4(6)(13);

	fa_4_0_14: fa
		port map(
			a => dadda_tree_4(0)(14),
			b => dadda_tree_4(1)(14),
			ci => dadda_tree_4(2)(14),
			s => dadda_tree_3(2)(14),
			co => dadda_tree_3(0)(15)
	);

	fa_4_3_14: fa
		port map(
			a => dadda_tree_4(3)(14),
			b => dadda_tree_4(4)(14),
			ci => dadda_tree_4(5)(14),
			s => dadda_tree_3(3)(14),
			co => dadda_tree_3(1)(15)
	);

	ha_4_6_14: ha
		port map(
			a => dadda_tree_4(6)(14),
			b => dadda_tree_4(7)(14),
			s => dadda_tree_3(4)(14),
			co => dadda_tree_3(2)(15)
	);

	dadda_tree_3(5)(14) <= dadda_tree_4(8)(14);

	fa_4_0_15: fa
		port map(
			a => dadda_tree_4(0)(15),
			b => dadda_tree_4(1)(15),
			ci => dadda_tree_4(2)(15),
			s => dadda_tree_3(3)(15),
			co => dadda_tree_3(0)(16)
	);

	fa_4_3_15: fa
		port map(
			a => dadda_tree_4(3)(15),
			b => dadda_tree_4(4)(15),
			ci => dadda_tree_4(5)(15),
			s => dadda_tree_3(4)(15),
			co => dadda_tree_3(1)(16)
	);

	ha_4_6_15: ha
		port map(
			a => dadda_tree_4(6)(15),
			b => dadda_tree_4(7)(15),
			s => dadda_tree_3(5)(15),
			co => dadda_tree_3(2)(16)
	);

	dadda_tree_3(0)(16) <= dadda_tree_4(0)(16);
	dadda_tree_3(0)(17) <= dadda_tree_4(0)(17);
	dadda_tree_3(1)(17) <= dadda_tree_4(1)(17);
	dadda_tree_3(0)(18) <= dadda_tree_4(0)(18);
	dadda_tree_3(1)(18) <= dadda_tree_4(1)(18);
	dadda_tree_3(2)(18) <= dadda_tree_4(2)(18);
	dadda_tree_3(0)(19) <= dadda_tree_4(0)(19);
	dadda_tree_3(1)(19) <= dadda_tree_4(1)(19);
	dadda_tree_3(2)(19) <= dadda_tree_4(2)(19);
	dadda_tree_3(3)(19) <= dadda_tree_4(3)(19);
	dadda_tree_3(0)(20) <= dadda_tree_4(0)(20);
	dadda_tree_3(1)(20) <= dadda_tree_4(1)(20);
	dadda_tree_3(2)(20) <= dadda_tree_4(2)(20);
	dadda_tree_3(3)(20) <= dadda_tree_4(3)(20);
	dadda_tree_3(4)(20) <= dadda_tree_4(4)(20);
	dadda_tree_3(0)(21) <= dadda_tree_4(0)(21);
	dadda_tree_3(1)(21) <= dadda_tree_4(1)(21);
	dadda_tree_3(2)(21) <= dadda_tree_4(2)(21);
	dadda_tree_3(3)(21) <= dadda_tree_4(3)(21);
	dadda_tree_3(4)(21) <= dadda_tree_4(4)(21);
	dadda_tree_3(5)(21) <= dadda_tree_4(5)(21);

	ha_4_0_22: ha
		port map(
			a => dadda_tree_4(0)(22),
			b => dadda_tree_4(1)(22),
			s => dadda_tree_3(0)(22),
			co => dadda_tree_3(0)(23)
	);

	dadda_tree_3(1)(22) <= dadda_tree_4(2)(22);
	dadda_tree_3(2)(22) <= dadda_tree_4(3)(22);
	dadda_tree_3(3)(22) <= dadda_tree_4(4)(22);
	dadda_tree_3(4)(22) <= dadda_tree_4(5)(22);
	dadda_tree_3(5)(22) <= dadda_tree_4(6)(22);

	fa_4_0_23: fa
		port map(
			a => dadda_tree_4(0)(23),
			b => dadda_tree_4(1)(23),
			ci => dadda_tree_4(2)(23),
			s => dadda_tree_3(1)(23),
			co => dadda_tree_3(0)(24)
	);

	ha_4_3_23: ha
		port map(
			a => dadda_tree_4(3)(23),
			b => dadda_tree_4(4)(23),
			s => dadda_tree_3(2)(23),
			co => dadda_tree_3(1)(24)
	);

	dadda_tree_3(3)(23) <= dadda_tree_4(5)(23);
	dadda_tree_3(4)(23) <= dadda_tree_4(6)(23);
	dadda_tree_3(5)(23) <= dadda_tree_4(7)(23);
	dadda_tree_3(0)(24) <= dadda_tree_4(0)(24);
	dadda_tree_3(0)(25) <= dadda_tree_4(0)(25);
	dadda_tree_3(1)(25) <= dadda_tree_4(1)(25);
	dadda_tree_3(0)(26) <= dadda_tree_4(0)(26);
	dadda_tree_3(1)(26) <= dadda_tree_4(1)(26);
	dadda_tree_3(2)(26) <= dadda_tree_4(2)(26);
	dadda_tree_3(0)(27) <= dadda_tree_4(0)(27);
	dadda_tree_3(1)(27) <= dadda_tree_4(1)(27);
	dadda_tree_3(2)(27) <= dadda_tree_4(2)(27);
	dadda_tree_3(3)(27) <= dadda_tree_4(3)(27);
	dadda_tree_3(0)(28) <= dadda_tree_4(0)(28);
	dadda_tree_3(1)(28) <= dadda_tree_4(1)(28);
	dadda_tree_3(2)(28) <= dadda_tree_4(2)(28);
	dadda_tree_3(3)(28) <= dadda_tree_4(3)(28);
	dadda_tree_3(4)(28) <= dadda_tree_4(4)(28);
	dadda_tree_3(0)(29) <= dadda_tree_4(0)(29);
	dadda_tree_3(1)(29) <= dadda_tree_4(1)(29);
	dadda_tree_3(2)(29) <= dadda_tree_4(2)(29);
	dadda_tree_3(3)(29) <= dadda_tree_4(3)(29);
	dadda_tree_3(4)(29) <= dadda_tree_4(4)(29);
	dadda_tree_3(5)(29) <= dadda_tree_4(5)(29);

	ha_4_0_30: ha
		port map(
			a => dadda_tree_4(0)(30),
			b => dadda_tree_4(1)(30),
			s => dadda_tree_3(0)(30),
			co => dadda_tree_3(0)(31)
	);

	dadda_tree_3(1)(30) <= dadda_tree_4(2)(30);
	dadda_tree_3(2)(30) <= dadda_tree_4(3)(30);
	dadda_tree_3(3)(30) <= dadda_tree_4(4)(30);
	dadda_tree_3(4)(30) <= dadda_tree_4(5)(30);
	dadda_tree_3(5)(30) <= dadda_tree_4(6)(30);

	fa_4_0_31: fa
		port map(
			a => dadda_tree_4(0)(31),
			b => dadda_tree_4(1)(31),
			ci => dadda_tree_4(2)(31),
			s => dadda_tree_3(1)(31),
			co => dadda_tree_3(0)(32)
	);

	ha_4_3_31: ha
		port map(
			a => dadda_tree_4(3)(31),
			b => dadda_tree_4(4)(31),
			s => dadda_tree_3(2)(31),
			co => dadda_tree_3(1)(32)
	);

	dadda_tree_3(3)(31) <= dadda_tree_4(5)(31);
	dadda_tree_3(4)(31) <= dadda_tree_4(6)(31);
	dadda_tree_3(5)(31) <= dadda_tree_4(7)(31);

	fa_4_0_32: fa
		port map(
			a => dadda_tree_4(0)(32),
			b => dadda_tree_4(1)(32),
			ci => dadda_tree_4(2)(32),
			s => dadda_tree_3(2)(32),
			co => dadda_tree_3(0)(33)
	);

	fa_4_3_32: fa
		port map(
			a => dadda_tree_4(3)(32),
			b => dadda_tree_4(4)(32),
			ci => dadda_tree_4(5)(32),
			s => dadda_tree_3(3)(32),
			co => dadda_tree_3(1)(33)
	);
	dadda_tree_3(4)(32) <= dadda_tree_4(6)(32);
	dadda_tree_3(5)(32) <= dadda_tree_4(7)(32);

	fa_4_0_33: fa
		port map(
			a => dadda_tree_4(0)(33),
			b => dadda_tree_4(1)(33),
			ci => dadda_tree_4(2)(33),
			s => dadda_tree_3(2)(33),
			co => dadda_tree_3(0)(34)
	);

	fa_4_3_33: fa
		port map(
			a => dadda_tree_4(3)(33),
			b => dadda_tree_4(4)(33),
			ci => dadda_tree_4(5)(33),
			s => dadda_tree_3(3)(33),
			co => dadda_tree_3(1)(34)
	);
	dadda_tree_3(4)(33) <= dadda_tree_4(6)(33);
	dadda_tree_3(5)(33) <= dadda_tree_4(7)(33);

	fa_4_0_34: fa
		port map(
			a => dadda_tree_4(0)(34),
			b => dadda_tree_4(1)(34),
			ci => dadda_tree_4(2)(34),
			s => dadda_tree_3(2)(34),
			co => dadda_tree_3(0)(35)
	);

	fa_4_3_34: fa
		port map(
			a => dadda_tree_4(3)(34),
			b => dadda_tree_4(4)(34),
			ci => dadda_tree_4(5)(34),
			s => dadda_tree_3(3)(34),
			co => dadda_tree_3(1)(35)
	);
	dadda_tree_3(4)(34) <= dadda_tree_4(6)(34);
	dadda_tree_3(5)(34) <= dadda_tree_4(7)(34);

	fa_4_0_35: fa
		port map(
			a => dadda_tree_4(0)(35),
			b => dadda_tree_4(1)(35),
			ci => dadda_tree_4(2)(35),
			s => dadda_tree_3(2)(35),
			co => dadda_tree_3(0)(36)
	);

	fa_4_3_35: fa
		port map(
			a => dadda_tree_4(3)(35),
			b => dadda_tree_4(4)(35),
			ci => dadda_tree_4(5)(35),
			s => dadda_tree_3(3)(35),
			co => dadda_tree_3(1)(36)
	);
	dadda_tree_3(4)(35) <= dadda_tree_4(6)(35);
	dadda_tree_3(5)(35) <= dadda_tree_4(7)(35);

	fa_4_0_36: fa
		port map(
			a => dadda_tree_4(0)(36),
			b => dadda_tree_4(1)(36),
			ci => dadda_tree_4(2)(36),
			s => dadda_tree_3(2)(36),
			co => dadda_tree_3(0)(37)
	);

	fa_4_3_36: fa
		port map(
			a => dadda_tree_4(3)(36),
			b => dadda_tree_4(4)(36),
			ci => dadda_tree_4(5)(36),
			s => dadda_tree_3(3)(36),
			co => dadda_tree_3(1)(37)
	);
	dadda_tree_3(4)(36) <= dadda_tree_4(6)(36);
	dadda_tree_3(5)(36) <= dadda_tree_4(7)(36);

	fa_4_0_37: fa
		port map(
			a => dadda_tree_4(0)(37),
			b => dadda_tree_4(1)(37),
			ci => dadda_tree_4(2)(37),
			s => dadda_tree_3(2)(37),
			co => dadda_tree_3(0)(38)
	);

	ha_4_3_37: ha
		port map(
			a => dadda_tree_4(3)(37),
			b => dadda_tree_4(4)(37),
			s => dadda_tree_3(3)(37),
			co => dadda_tree_3(1)(38)
	);

	dadda_tree_3(4)(37) <= dadda_tree_4(5)(37);
	dadda_tree_3(5)(37) <= dadda_tree_4(6)(37);

	fa_4_0_38: fa
		port map(
			a => dadda_tree_4(0)(38),
			b => dadda_tree_4(1)(38),
			ci => dadda_tree_4(2)(38),
			s => dadda_tree_3(2)(38),
			co => dadda_tree_3(0)(39)
	);
	dadda_tree_3(3)(38) <= dadda_tree_4(3)(38);
	dadda_tree_3(4)(38) <= dadda_tree_4(4)(38);
	dadda_tree_3(5)(38) <= dadda_tree_4(5)(38);
	dadda_tree_3(0)(39) <= dadda_tree_4(0)(39);
	dadda_tree_3(1)(39) <= dadda_tree_4(1)(39);
	dadda_tree_3(2)(39) <= dadda_tree_4(2)(39);
	dadda_tree_3(3)(39) <= dadda_tree_4(3)(39);
	dadda_tree_3(4)(39) <= dadda_tree_4(4)(39);
	dadda_tree_3(0)(40) <= dadda_tree_4(0)(40);
	dadda_tree_3(1)(40) <= dadda_tree_4(1)(40);
	dadda_tree_3(2)(40) <= dadda_tree_4(2)(40);
	dadda_tree_3(3)(40) <= dadda_tree_4(3)(40);
	dadda_tree_3(0)(41) <= dadda_tree_4(0)(41);
	dadda_tree_3(1)(41) <= dadda_tree_4(1)(41);
	dadda_tree_3(2)(41) <= dadda_tree_4(2)(41);
	dadda_tree_3(0)(42) <= dadda_tree_4(0)(42);
	dadda_tree_3(1)(42) <= dadda_tree_4(1)(42);
	dadda_tree_3(0)(43) <= dadda_tree_4(0)(43);
	dadda_tree_3(1)(43) <= dadda_tree_4(1)(43);
	dadda_tree_3(0)(44) <= dadda_tree_4(0)(44);
	dadda_tree_3(1)(44) <= dadda_tree_4(1)(44);
	dadda_tree_3(2)(44) <= dadda_tree_4(2)(44);
	dadda_tree_3(3)(44) <= dadda_tree_4(3)(44);
	dadda_tree_3(4)(44) <= dadda_tree_4(4)(44);
	dadda_tree_3(0)(45) <= dadda_tree_4(0)(45);
	dadda_tree_3(1)(45) <= dadda_tree_4(1)(45);
	dadda_tree_3(2)(45) <= dadda_tree_4(2)(45);
	dadda_tree_3(3)(45) <= dadda_tree_4(3)(45);
	dadda_tree_3(4)(45) <= dadda_tree_4(4)(45);
	dadda_tree_3(5)(45) <= dadda_tree_4(5)(45);
	dadda_tree_3(0)(46) <= dadda_tree_4(0)(46);
	dadda_tree_3(1)(46) <= dadda_tree_4(1)(46);
	dadda_tree_3(2)(46) <= dadda_tree_4(2)(46);
	dadda_tree_3(3)(46) <= dadda_tree_4(3)(46);
	dadda_tree_3(4)(46) <= dadda_tree_4(4)(46);
	dadda_tree_3(5)(46) <= dadda_tree_4(5)(46);
	dadda_tree_3(0)(47) <= dadda_tree_4(0)(47);
	dadda_tree_3(1)(47) <= dadda_tree_4(1)(47);
	dadda_tree_3(2)(47) <= dadda_tree_4(2)(47);
	dadda_tree_3(3)(47) <= dadda_tree_4(3)(47);
	dadda_tree_3(4)(47) <= dadda_tree_4(4)(47);
	dadda_tree_3(0)(48) <= dadda_tree_4(0)(48);
	dadda_tree_3(1)(48) <= dadda_tree_4(1)(48);
	dadda_tree_3(2)(48) <= dadda_tree_4(2)(48);
	dadda_tree_3(3)(48) <= dadda_tree_4(3)(48);
	dadda_tree_3(0)(49) <= dadda_tree_4(0)(49);
	dadda_tree_3(1)(49) <= dadda_tree_4(1)(49);
	dadda_tree_3(2)(49) <= dadda_tree_4(2)(49);
	dadda_tree_3(0)(50) <= dadda_tree_4(0)(50);
	dadda_tree_3(1)(50) <= dadda_tree_4(1)(50);

	fa_4_0_51: fa
		port map(
			a => dadda_tree_4(0)(51),
			b => dadda_tree_4(1)(51),
			ci => dadda_tree_4(2)(51),
			s => dadda_tree_3(0)(51),
			co => dadda_tree_3(0)(52)
	);
	dadda_tree_3(1)(51) <= dadda_tree_4(3)(51);
	dadda_tree_3(2)(51) <= dadda_tree_4(4)(51);
	dadda_tree_3(3)(51) <= dadda_tree_4(5)(51);
	dadda_tree_3(4)(51) <= dadda_tree_4(6)(51);
	dadda_tree_3(5)(51) <= dadda_tree_4(7)(51);

	fa_4_0_52: fa
		port map(
			a => dadda_tree_4(0)(52),
			b => dadda_tree_4(1)(52),
			ci => dadda_tree_4(2)(52),
			s => dadda_tree_3(1)(52),
			co => dadda_tree_3(0)(53)
	);

	ha_4_3_52: ha
		port map(
			a => dadda_tree_4(3)(52),
			b => dadda_tree_4(4)(52),
			s => dadda_tree_3(2)(52),
			co => dadda_tree_3(1)(53)
	);

	dadda_tree_3(3)(52) <= dadda_tree_4(5)(52);
	dadda_tree_3(4)(52) <= dadda_tree_4(6)(52);
	dadda_tree_3(5)(52) <= dadda_tree_4(7)(52);

	fa_4_0_53: fa
		port map(
			a => dadda_tree_4(0)(53),
			b => dadda_tree_4(1)(53),
			ci => dadda_tree_4(2)(53),
			s => dadda_tree_3(2)(53),
			co => dadda_tree_3(0)(54)
	);

	ha_4_3_53: ha
		port map(
			a => dadda_tree_4(3)(53),
			b => dadda_tree_4(4)(53),
			s => dadda_tree_3(3)(53),
			co => dadda_tree_3(1)(54)
	);

	dadda_tree_3(4)(53) <= dadda_tree_4(5)(53);
	dadda_tree_3(5)(53) <= dadda_tree_4(6)(53);

	fa_4_0_54: fa
		port map(
			a => dadda_tree_4(0)(54),
			b => dadda_tree_4(1)(54),
			ci => dadda_tree_4(2)(54),
			s => dadda_tree_3(2)(54),
			co => dadda_tree_3(0)(55)
	);

	ha_4_3_54: ha
		port map(
			a => dadda_tree_4(3)(54),
			b => dadda_tree_4(4)(54),
			s => dadda_tree_3(3)(54),
			co => dadda_tree_3(1)(55)
	);

	dadda_tree_3(4)(54) <= dadda_tree_4(5)(54);
	dadda_tree_3(5)(54) <= dadda_tree_4(6)(54);

	fa_4_0_55: fa
		port map(
			a => dadda_tree_4(0)(55),
			b => dadda_tree_4(1)(55),
			ci => dadda_tree_4(2)(55),
			s => dadda_tree_3(2)(55),
			co => dadda_tree_3(0)(56)
	);
	dadda_tree_3(3)(55) <= dadda_tree_4(3)(55);
	dadda_tree_3(4)(55) <= dadda_tree_4(4)(55);
	dadda_tree_3(5)(55) <= dadda_tree_4(5)(55);

	ha_4_0_56: ha
		port map(
			a => dadda_tree_4(0)(56),
			b => dadda_tree_4(1)(56),
			s => dadda_tree_3(1)(56),
			co => dadda_tree_3(0)(57)
	);

	dadda_tree_3(2)(56) <= dadda_tree_4(2)(56);
	dadda_tree_3(3)(56) <= dadda_tree_4(3)(56);
	dadda_tree_3(4)(56) <= dadda_tree_4(4)(56);
	dadda_tree_3(5)(56) <= dadda_tree_4(5)(56);
	dadda_tree_3(0)(57) <= dadda_tree_4(0)(57);
	dadda_tree_3(1)(57) <= dadda_tree_4(1)(57);
	dadda_tree_3(2)(57) <= dadda_tree_4(2)(57);
	dadda_tree_3(3)(57) <= dadda_tree_4(3)(57);
	dadda_tree_3(4)(57) <= dadda_tree_4(4)(57);
	dadda_tree_3(0)(58) <= dadda_tree_4(0)(58);
	dadda_tree_3(1)(58) <= dadda_tree_4(1)(58);
	dadda_tree_3(2)(58) <= dadda_tree_4(2)(58);
	dadda_tree_3(3)(58) <= dadda_tree_4(3)(58);
	dadda_tree_3(4)(58) <= dadda_tree_4(4)(58);
	dadda_tree_3(0)(59) <= dadda_tree_4(0)(59);
	dadda_tree_3(1)(59) <= dadda_tree_4(1)(59);
	dadda_tree_3(2)(59) <= dadda_tree_4(2)(59);
	dadda_tree_3(3)(59) <= dadda_tree_4(3)(59);
	dadda_tree_3(0)(60) <= dadda_tree_4(0)(60);
	dadda_tree_3(1)(60) <= dadda_tree_4(1)(60);
	dadda_tree_3(2)(60) <= dadda_tree_4(2)(60);
	dadda_tree_3(3)(60) <= dadda_tree_4(3)(60);
	dadda_tree_3(0)(61) <= dadda_tree_4(0)(61);
	dadda_tree_3(1)(61) <= dadda_tree_4(1)(61);
	dadda_tree_3(2)(61) <= dadda_tree_4(2)(61);
	dadda_tree_3(0)(62) <= dadda_tree_4(0)(62);
	dadda_tree_3(1)(62) <= dadda_tree_4(1)(62);
	dadda_tree_3(2)(62) <= dadda_tree_4(2)(62);
	dadda_tree_3(0)(63) <= dadda_tree_4(0)(63);
	dadda_tree_3(1)(63) <= dadda_tree_4(1)(63);
	dadda_tree_2(0)(0) <= dadda_tree_3(0)(0);
	dadda_tree_2(1)(0) <= dadda_tree_3(1)(0);
	dadda_tree_2(0)(1) <= dadda_tree_3(0)(1);
	dadda_tree_2(0)(2) <= dadda_tree_3(0)(2);
	dadda_tree_2(1)(2) <= dadda_tree_3(1)(2);
	dadda_tree_2(2)(2) <= dadda_tree_3(2)(2);
	dadda_tree_2(0)(3) <= dadda_tree_3(0)(3);
	dadda_tree_2(1)(3) <= dadda_tree_3(1)(3);
	dadda_tree_2(0)(4) <= dadda_tree_3(0)(4);
	dadda_tree_2(1)(4) <= dadda_tree_3(1)(4);
	dadda_tree_2(2)(4) <= dadda_tree_3(2)(4);
	dadda_tree_2(3)(4) <= dadda_tree_3(3)(4);
	dadda_tree_2(0)(5) <= dadda_tree_3(0)(5);
	dadda_tree_2(1)(5) <= dadda_tree_3(1)(5);
	dadda_tree_2(2)(5) <= dadda_tree_3(2)(5);

	ha_3_0_6: ha
		port map(
			a => dadda_tree_3(0)(6),
			b => dadda_tree_3(1)(6),
			s => dadda_tree_2(0)(6),
			co => dadda_tree_2(0)(7)
	);

	dadda_tree_2(1)(6) <= dadda_tree_3(2)(6);
	dadda_tree_2(2)(6) <= dadda_tree_3(3)(6);
	dadda_tree_2(3)(6) <= dadda_tree_3(4)(6);

	ha_3_0_7: ha
		port map(
			a => dadda_tree_3(0)(7),
			b => dadda_tree_3(1)(7),
			s => dadda_tree_2(1)(7),
			co => dadda_tree_2(0)(8)
	);

	dadda_tree_2(2)(7) <= dadda_tree_3(2)(7);
	dadda_tree_2(3)(7) <= dadda_tree_3(3)(7);

	fa_3_0_8: fa
		port map(
			a => dadda_tree_3(0)(8),
			b => dadda_tree_3(1)(8),
			ci => dadda_tree_3(2)(8),
			s => dadda_tree_2(1)(8),
			co => dadda_tree_2(0)(9)
	);

	ha_3_3_8: ha
		port map(
			a => dadda_tree_3(3)(8),
			b => dadda_tree_3(4)(8),
			s => dadda_tree_2(2)(8),
			co => dadda_tree_2(1)(9)
	);

	dadda_tree_2(3)(8) <= dadda_tree_3(5)(8);

	fa_3_0_9: fa
		port map(
			a => dadda_tree_3(0)(9),
			b => dadda_tree_3(1)(9),
			ci => dadda_tree_3(2)(9),
			s => dadda_tree_2(2)(9),
			co => dadda_tree_2(0)(10)
	);

	ha_3_3_9: ha
		port map(
			a => dadda_tree_3(3)(9),
			b => dadda_tree_3(4)(9),
			s => dadda_tree_2(3)(9),
			co => dadda_tree_2(1)(10)
	);

	dadda_tree_2(0)(10) <= dadda_tree_3(0)(10);
	dadda_tree_2(0)(11) <= dadda_tree_3(0)(11);
	dadda_tree_2(1)(11) <= dadda_tree_3(1)(11);
	dadda_tree_2(0)(12) <= dadda_tree_3(0)(12);
	dadda_tree_2(1)(12) <= dadda_tree_3(1)(12);
	dadda_tree_2(2)(12) <= dadda_tree_3(2)(12);
	dadda_tree_2(0)(13) <= dadda_tree_3(0)(13);
	dadda_tree_2(1)(13) <= dadda_tree_3(1)(13);
	dadda_tree_2(2)(13) <= dadda_tree_3(2)(13);
	dadda_tree_2(3)(13) <= dadda_tree_3(3)(13);

	ha_3_0_14: ha
		port map(
			a => dadda_tree_3(0)(14),
			b => dadda_tree_3(1)(14),
			s => dadda_tree_2(0)(14),
			co => dadda_tree_2(0)(15)
	);

	dadda_tree_2(1)(14) <= dadda_tree_3(2)(14);
	dadda_tree_2(2)(14) <= dadda_tree_3(3)(14);
	dadda_tree_2(3)(14) <= dadda_tree_3(4)(14);

	fa_3_0_15: fa
		port map(
			a => dadda_tree_3(0)(15),
			b => dadda_tree_3(1)(15),
			ci => dadda_tree_3(2)(15),
			s => dadda_tree_2(1)(15),
			co => dadda_tree_2(0)(16)
	);

	ha_3_3_15: ha
		port map(
			a => dadda_tree_3(3)(15),
			b => dadda_tree_3(4)(15),
			s => dadda_tree_2(2)(15),
			co => dadda_tree_2(1)(16)
	);

	dadda_tree_2(3)(15) <= dadda_tree_3(5)(15);
	dadda_tree_2(0)(16) <= dadda_tree_3(0)(16);
	dadda_tree_2(0)(17) <= dadda_tree_3(0)(17);
	dadda_tree_2(1)(17) <= dadda_tree_3(1)(17);
	dadda_tree_2(0)(18) <= dadda_tree_3(0)(18);
	dadda_tree_2(1)(18) <= dadda_tree_3(1)(18);
	dadda_tree_2(2)(18) <= dadda_tree_3(2)(18);
	dadda_tree_2(0)(19) <= dadda_tree_3(0)(19);
	dadda_tree_2(1)(19) <= dadda_tree_3(1)(19);
	dadda_tree_2(2)(19) <= dadda_tree_3(2)(19);
	dadda_tree_2(3)(19) <= dadda_tree_3(3)(19);

	ha_3_0_20: ha
		port map(
			a => dadda_tree_3(0)(20),
			b => dadda_tree_3(1)(20),
			s => dadda_tree_2(0)(20),
			co => dadda_tree_2(0)(21)
	);

	dadda_tree_2(1)(20) <= dadda_tree_3(2)(20);
	dadda_tree_2(2)(20) <= dadda_tree_3(3)(20);
	dadda_tree_2(3)(20) <= dadda_tree_3(4)(20);

	fa_3_0_21: fa
		port map(
			a => dadda_tree_3(0)(21),
			b => dadda_tree_3(1)(21),
			ci => dadda_tree_3(2)(21),
			s => dadda_tree_2(1)(21),
			co => dadda_tree_2(0)(22)
	);

	ha_3_3_21: ha
		port map(
			a => dadda_tree_3(3)(21),
			b => dadda_tree_3(4)(21),
			s => dadda_tree_2(2)(21),
			co => dadda_tree_2(1)(22)
	);

	dadda_tree_2(3)(21) <= dadda_tree_3(5)(21);
	dadda_tree_2(0)(22) <= dadda_tree_3(0)(22);
	dadda_tree_2(0)(23) <= dadda_tree_3(0)(23);
	dadda_tree_2(1)(23) <= dadda_tree_3(1)(23);
	dadda_tree_2(2)(23) <= dadda_tree_3(2)(23);
	dadda_tree_2(0)(24) <= dadda_tree_3(0)(24);
	dadda_tree_2(0)(25) <= dadda_tree_3(0)(25);
	dadda_tree_2(1)(25) <= dadda_tree_3(1)(25);
	dadda_tree_2(0)(26) <= dadda_tree_3(0)(26);
	dadda_tree_2(1)(26) <= dadda_tree_3(1)(26);
	dadda_tree_2(2)(26) <= dadda_tree_3(2)(26);
	dadda_tree_2(0)(27) <= dadda_tree_3(0)(27);
	dadda_tree_2(1)(27) <= dadda_tree_3(1)(27);
	dadda_tree_2(2)(27) <= dadda_tree_3(2)(27);
	dadda_tree_2(3)(27) <= dadda_tree_3(3)(27);

	ha_3_0_28: ha
		port map(
			a => dadda_tree_3(0)(28),
			b => dadda_tree_3(1)(28),
			s => dadda_tree_2(0)(28),
			co => dadda_tree_2(0)(29)
	);

	dadda_tree_2(1)(28) <= dadda_tree_3(2)(28);
	dadda_tree_2(2)(28) <= dadda_tree_3(3)(28);
	dadda_tree_2(3)(28) <= dadda_tree_3(4)(28);

	fa_3_0_29: fa
		port map(
			a => dadda_tree_3(0)(29),
			b => dadda_tree_3(1)(29),
			ci => dadda_tree_3(2)(29),
			s => dadda_tree_2(1)(29),
			co => dadda_tree_2(0)(30)
	);

	ha_3_3_29: ha
		port map(
			a => dadda_tree_3(3)(29),
			b => dadda_tree_3(4)(29),
			s => dadda_tree_2(2)(29),
			co => dadda_tree_2(1)(30)
	);

	dadda_tree_2(3)(29) <= dadda_tree_3(5)(29);
	dadda_tree_2(0)(30) <= dadda_tree_3(0)(30);
	dadda_tree_2(0)(31) <= dadda_tree_3(0)(31);
	dadda_tree_2(1)(31) <= dadda_tree_3(1)(31);
	dadda_tree_2(2)(31) <= dadda_tree_3(2)(31);
	dadda_tree_2(0)(32) <= dadda_tree_3(0)(32);
	dadda_tree_2(1)(32) <= dadda_tree_3(1)(32);
	dadda_tree_2(2)(32) <= dadda_tree_3(2)(32);
	dadda_tree_2(3)(32) <= dadda_tree_3(3)(32);
	dadda_tree_2(0)(33) <= dadda_tree_3(0)(33);
	dadda_tree_2(1)(33) <= dadda_tree_3(1)(33);
	dadda_tree_2(2)(33) <= dadda_tree_3(2)(33);
	dadda_tree_2(3)(33) <= dadda_tree_3(3)(33);
	dadda_tree_2(0)(34) <= dadda_tree_3(0)(34);
	dadda_tree_2(1)(34) <= dadda_tree_3(1)(34);
	dadda_tree_2(2)(34) <= dadda_tree_3(2)(34);
	dadda_tree_2(3)(34) <= dadda_tree_3(3)(34);
	dadda_tree_2(0)(35) <= dadda_tree_3(0)(35);
	dadda_tree_2(1)(35) <= dadda_tree_3(1)(35);
	dadda_tree_2(2)(35) <= dadda_tree_3(2)(35);
	dadda_tree_2(3)(35) <= dadda_tree_3(3)(35);
	dadda_tree_2(0)(36) <= dadda_tree_3(0)(36);
	dadda_tree_2(1)(36) <= dadda_tree_3(1)(36);
	dadda_tree_2(2)(36) <= dadda_tree_3(2)(36);
	dadda_tree_2(3)(36) <= dadda_tree_3(3)(36);
	dadda_tree_2(0)(37) <= dadda_tree_3(0)(37);
	dadda_tree_2(1)(37) <= dadda_tree_3(1)(37);
	dadda_tree_2(2)(37) <= dadda_tree_3(2)(37);
	dadda_tree_2(3)(37) <= dadda_tree_3(3)(37);
	dadda_tree_2(0)(38) <= dadda_tree_3(0)(38);
	dadda_tree_2(1)(38) <= dadda_tree_3(1)(38);
	dadda_tree_2(2)(38) <= dadda_tree_3(2)(38);

	ha_3_0_39: ha
		port map(
			a => dadda_tree_3(0)(39),
			b => dadda_tree_3(1)(39),
			s => dadda_tree_2(0)(39),
			co => dadda_tree_2(0)(40)
	);

	dadda_tree_2(1)(39) <= dadda_tree_3(2)(39);
	dadda_tree_2(2)(39) <= dadda_tree_3(3)(39);
	dadda_tree_2(3)(39) <= dadda_tree_3(4)(39);

	ha_3_0_40: ha
		port map(
			a => dadda_tree_3(0)(40),
			b => dadda_tree_3(1)(40),
			s => dadda_tree_2(1)(40),
			co => dadda_tree_2(0)(41)
	);

	dadda_tree_2(2)(40) <= dadda_tree_3(2)(40);
	dadda_tree_2(3)(40) <= dadda_tree_3(3)(40);
	dadda_tree_2(0)(41) <= dadda_tree_3(0)(41);
	dadda_tree_2(1)(41) <= dadda_tree_3(1)(41);
	dadda_tree_2(2)(41) <= dadda_tree_3(2)(41);
	dadda_tree_2(0)(42) <= dadda_tree_3(0)(42);
	dadda_tree_2(1)(42) <= dadda_tree_3(1)(42);
	dadda_tree_2(0)(43) <= dadda_tree_3(0)(43);
	dadda_tree_2(1)(43) <= dadda_tree_3(1)(43);

	ha_3_0_44: ha
		port map(
			a => dadda_tree_3(0)(44),
			b => dadda_tree_3(1)(44),
			s => dadda_tree_2(0)(44),
			co => dadda_tree_2(0)(45)
	);

	dadda_tree_2(1)(44) <= dadda_tree_3(2)(44);
	dadda_tree_2(2)(44) <= dadda_tree_3(3)(44);
	dadda_tree_2(3)(44) <= dadda_tree_3(4)(44);

	fa_3_0_45: fa
		port map(
			a => dadda_tree_3(0)(45),
			b => dadda_tree_3(1)(45),
			ci => dadda_tree_3(2)(45),
			s => dadda_tree_2(1)(45),
			co => dadda_tree_2(0)(46)
	);

	ha_3_3_45: ha
		port map(
			a => dadda_tree_3(3)(45),
			b => dadda_tree_3(4)(45),
			s => dadda_tree_2(2)(45),
			co => dadda_tree_2(1)(46)
	);

	dadda_tree_2(3)(45) <= dadda_tree_3(5)(45);

	fa_3_0_46: fa
		port map(
			a => dadda_tree_3(0)(46),
			b => dadda_tree_3(1)(46),
			ci => dadda_tree_3(2)(46),
			s => dadda_tree_2(2)(46),
			co => dadda_tree_2(0)(47)
	);

	fa_3_3_46: fa
		port map(
			a => dadda_tree_3(3)(46),
			b => dadda_tree_3(4)(46),
			ci => dadda_tree_3(5)(46),
			s => dadda_tree_2(3)(46),
			co => dadda_tree_2(1)(47)
	);

	fa_3_0_47: fa
		port map(
			a => dadda_tree_3(0)(47),
			b => dadda_tree_3(1)(47),
			ci => dadda_tree_3(2)(47),
			s => dadda_tree_2(2)(47),
			co => dadda_tree_2(0)(48)
	);

	ha_3_3_47: ha
		port map(
			a => dadda_tree_3(3)(47),
			b => dadda_tree_3(4)(47),
			s => dadda_tree_2(3)(47),
			co => dadda_tree_2(1)(48)
	);


	fa_3_0_48: fa
		port map(
			a => dadda_tree_3(0)(48),
			b => dadda_tree_3(1)(48),
			ci => dadda_tree_3(2)(48),
			s => dadda_tree_2(2)(48),
			co => dadda_tree_2(0)(49)
	);
	dadda_tree_2(3)(48) <= dadda_tree_3(3)(48);
	dadda_tree_2(0)(49) <= dadda_tree_3(0)(49);
	dadda_tree_2(1)(49) <= dadda_tree_3(1)(49);
	dadda_tree_2(2)(49) <= dadda_tree_3(2)(49);
	dadda_tree_2(0)(50) <= dadda_tree_3(0)(50);
	dadda_tree_2(1)(50) <= dadda_tree_3(1)(50);
	dadda_tree_2(0)(51) <= dadda_tree_3(0)(51);
	dadda_tree_2(0)(52) <= dadda_tree_3(0)(52);
	dadda_tree_2(1)(52) <= dadda_tree_3(1)(52);
	dadda_tree_2(2)(52) <= dadda_tree_3(2)(52);
	dadda_tree_2(0)(53) <= dadda_tree_3(0)(53);
	dadda_tree_2(1)(53) <= dadda_tree_3(1)(53);
	dadda_tree_2(2)(53) <= dadda_tree_3(2)(53);
	dadda_tree_2(3)(53) <= dadda_tree_3(3)(53);
	dadda_tree_2(0)(54) <= dadda_tree_3(0)(54);
	dadda_tree_2(1)(54) <= dadda_tree_3(1)(54);
	dadda_tree_2(2)(54) <= dadda_tree_3(2)(54);
	dadda_tree_2(3)(54) <= dadda_tree_3(3)(54);
	dadda_tree_2(0)(55) <= dadda_tree_3(0)(55);
	dadda_tree_2(1)(55) <= dadda_tree_3(1)(55);
	dadda_tree_2(2)(55) <= dadda_tree_3(2)(55);
	dadda_tree_2(0)(56) <= dadda_tree_3(0)(56);
	dadda_tree_2(1)(56) <= dadda_tree_3(1)(56);

	ha_3_0_57: ha
		port map(
			a => dadda_tree_3(0)(57),
			b => dadda_tree_3(1)(57),
			s => dadda_tree_2(0)(57),
			co => dadda_tree_2(0)(58)
	);

	dadda_tree_2(1)(57) <= dadda_tree_3(2)(57);
	dadda_tree_2(2)(57) <= dadda_tree_3(3)(57);
	dadda_tree_2(3)(57) <= dadda_tree_3(4)(57);

	fa_3_0_58: fa
		port map(
			a => dadda_tree_3(0)(58),
			b => dadda_tree_3(1)(58),
			ci => dadda_tree_3(2)(58),
			s => dadda_tree_2(1)(58),
			co => dadda_tree_2(0)(59)
	);
	dadda_tree_2(2)(58) <= dadda_tree_3(3)(58);
	dadda_tree_2(3)(58) <= dadda_tree_3(4)(58);

	ha_3_0_59: ha
		port map(
			a => dadda_tree_3(0)(59),
			b => dadda_tree_3(1)(59),
			s => dadda_tree_2(1)(59),
			co => dadda_tree_2(0)(60)
	);

	dadda_tree_2(2)(59) <= dadda_tree_3(2)(59);
	dadda_tree_2(3)(59) <= dadda_tree_3(3)(59);

	ha_3_0_60: ha
		port map(
			a => dadda_tree_3(0)(60),
			b => dadda_tree_3(1)(60),
			s => dadda_tree_2(1)(60),
			co => dadda_tree_2(0)(61)
	);

	dadda_tree_2(2)(60) <= dadda_tree_3(2)(60);
	dadda_tree_2(3)(60) <= dadda_tree_3(3)(60);
	dadda_tree_2(0)(61) <= dadda_tree_3(0)(61);
	dadda_tree_2(1)(61) <= dadda_tree_3(1)(61);
	dadda_tree_2(2)(61) <= dadda_tree_3(2)(61);
	dadda_tree_2(0)(62) <= dadda_tree_3(0)(62);
	dadda_tree_2(1)(62) <= dadda_tree_3(1)(62);
	dadda_tree_2(2)(62) <= dadda_tree_3(2)(62);
	dadda_tree_2(0)(63) <= dadda_tree_3(0)(63);
	dadda_tree_2(1)(63) <= dadda_tree_3(1)(63);
	dadda_tree_1(0)(0) <= dadda_tree_2(0)(0);
	dadda_tree_1(1)(0) <= dadda_tree_2(1)(0);
	dadda_tree_1(0)(1) <= dadda_tree_2(0)(1);
	dadda_tree_1(0)(2) <= dadda_tree_2(0)(2);
	dadda_tree_1(1)(2) <= dadda_tree_2(1)(2);
	dadda_tree_1(2)(2) <= dadda_tree_2(2)(2);
	dadda_tree_1(0)(3) <= dadda_tree_2(0)(3);
	dadda_tree_1(1)(3) <= dadda_tree_2(1)(3);

	ha_2_0_4: ha
		port map(
			a => dadda_tree_2(0)(4),
			b => dadda_tree_2(1)(4),
			s => dadda_tree_1(0)(4),
			co => dadda_tree_1(0)(5)
	);

	dadda_tree_1(1)(4) <= dadda_tree_2(2)(4);
	dadda_tree_1(2)(4) <= dadda_tree_2(3)(4);

	ha_2_0_5: ha
		port map(
			a => dadda_tree_2(0)(5),
			b => dadda_tree_2(1)(5),
			s => dadda_tree_1(1)(5),
			co => dadda_tree_1(0)(6)
	);

	dadda_tree_1(2)(5) <= dadda_tree_2(2)(5);
	dadda_tree_1(0)(6) <= dadda_tree_2(0)(6);
	dadda_tree_1(0)(7) <= dadda_tree_2(0)(7);
	dadda_tree_1(1)(7) <= dadda_tree_2(1)(7);
	dadda_tree_1(0)(8) <= dadda_tree_2(0)(8);
	dadda_tree_1(1)(8) <= dadda_tree_2(1)(8);
	dadda_tree_1(2)(8) <= dadda_tree_2(2)(8);

	ha_2_0_9: ha
		port map(
			a => dadda_tree_2(0)(9),
			b => dadda_tree_2(1)(9),
			s => dadda_tree_1(0)(9),
			co => dadda_tree_1(0)(10)
	);

	dadda_tree_1(1)(9) <= dadda_tree_2(2)(9);
	dadda_tree_1(2)(9) <= dadda_tree_2(3)(9);
	dadda_tree_1(0)(10) <= dadda_tree_2(0)(10);
	dadda_tree_1(0)(11) <= dadda_tree_2(0)(11);
	dadda_tree_1(1)(11) <= dadda_tree_2(1)(11);
	dadda_tree_1(0)(12) <= dadda_tree_2(0)(12);
	dadda_tree_1(1)(12) <= dadda_tree_2(1)(12);
	dadda_tree_1(2)(12) <= dadda_tree_2(2)(12);

	ha_2_0_13: ha
		port map(
			a => dadda_tree_2(0)(13),
			b => dadda_tree_2(1)(13),
			s => dadda_tree_1(0)(13),
			co => dadda_tree_1(0)(14)
	);

	dadda_tree_1(1)(13) <= dadda_tree_2(2)(13);
	dadda_tree_1(2)(13) <= dadda_tree_2(3)(13);
	dadda_tree_1(0)(14) <= dadda_tree_2(0)(14);
	dadda_tree_1(0)(15) <= dadda_tree_2(0)(15);
	dadda_tree_1(1)(15) <= dadda_tree_2(1)(15);
	dadda_tree_1(2)(15) <= dadda_tree_2(2)(15);
	dadda_tree_1(0)(16) <= dadda_tree_2(0)(16);
	dadda_tree_1(0)(17) <= dadda_tree_2(0)(17);
	dadda_tree_1(1)(17) <= dadda_tree_2(1)(17);
	dadda_tree_1(0)(18) <= dadda_tree_2(0)(18);
	dadda_tree_1(1)(18) <= dadda_tree_2(1)(18);
	dadda_tree_1(2)(18) <= dadda_tree_2(2)(18);

	ha_2_0_19: ha
		port map(
			a => dadda_tree_2(0)(19),
			b => dadda_tree_2(1)(19),
			s => dadda_tree_1(0)(19),
			co => dadda_tree_1(0)(20)
	);

	dadda_tree_1(1)(19) <= dadda_tree_2(2)(19);
	dadda_tree_1(2)(19) <= dadda_tree_2(3)(19);
	dadda_tree_1(0)(20) <= dadda_tree_2(0)(20);
	dadda_tree_1(0)(21) <= dadda_tree_2(0)(21);
	dadda_tree_1(1)(21) <= dadda_tree_2(1)(21);
	dadda_tree_1(2)(21) <= dadda_tree_2(2)(21);
	dadda_tree_1(0)(22) <= dadda_tree_2(0)(22);
	dadda_tree_1(0)(23) <= dadda_tree_2(0)(23);
	dadda_tree_1(1)(23) <= dadda_tree_2(1)(23);
	dadda_tree_1(2)(23) <= dadda_tree_2(2)(23);
	dadda_tree_1(0)(24) <= dadda_tree_2(0)(24);
	dadda_tree_1(0)(25) <= dadda_tree_2(0)(25);
	dadda_tree_1(1)(25) <= dadda_tree_2(1)(25);
	dadda_tree_1(0)(26) <= dadda_tree_2(0)(26);
	dadda_tree_1(1)(26) <= dadda_tree_2(1)(26);
	dadda_tree_1(2)(26) <= dadda_tree_2(2)(26);

	ha_2_0_27: ha
		port map(
			a => dadda_tree_2(0)(27),
			b => dadda_tree_2(1)(27),
			s => dadda_tree_1(0)(27),
			co => dadda_tree_1(0)(28)
	);

	dadda_tree_1(1)(27) <= dadda_tree_2(2)(27);
	dadda_tree_1(2)(27) <= dadda_tree_2(3)(27);
	dadda_tree_1(0)(28) <= dadda_tree_2(0)(28);
	dadda_tree_1(0)(29) <= dadda_tree_2(0)(29);
	dadda_tree_1(1)(29) <= dadda_tree_2(1)(29);
	dadda_tree_1(2)(29) <= dadda_tree_2(2)(29);
	dadda_tree_1(0)(30) <= dadda_tree_2(0)(30);
	dadda_tree_1(0)(31) <= dadda_tree_2(0)(31);
	dadda_tree_1(1)(31) <= dadda_tree_2(1)(31);
	dadda_tree_1(2)(31) <= dadda_tree_2(2)(31);

	ha_2_0_32: ha
		port map(
			a => dadda_tree_2(0)(32),
			b => dadda_tree_2(1)(32),
			s => dadda_tree_1(0)(32),
			co => dadda_tree_1(0)(33)
	);

	dadda_tree_1(1)(32) <= dadda_tree_2(2)(32);
	dadda_tree_1(2)(32) <= dadda_tree_2(3)(32);

	fa_2_0_33: fa
		port map(
			a => dadda_tree_2(0)(33),
			b => dadda_tree_2(1)(33),
			ci => dadda_tree_2(2)(33),
			s => dadda_tree_1(1)(33),
			co => dadda_tree_1(0)(34)
	);
	dadda_tree_1(2)(33) <= dadda_tree_2(3)(33);

	fa_2_0_34: fa
		port map(
			a => dadda_tree_2(0)(34),
			b => dadda_tree_2(1)(34),
			ci => dadda_tree_2(2)(34),
			s => dadda_tree_1(1)(34),
			co => dadda_tree_1(0)(35)
	);
	dadda_tree_1(2)(34) <= dadda_tree_2(3)(34);

	fa_2_0_35: fa
		port map(
			a => dadda_tree_2(0)(35),
			b => dadda_tree_2(1)(35),
			ci => dadda_tree_2(2)(35),
			s => dadda_tree_1(1)(35),
			co => dadda_tree_1(0)(36)
	);
	dadda_tree_1(2)(35) <= dadda_tree_2(3)(35);

	fa_2_0_36: fa
		port map(
			a => dadda_tree_2(0)(36),
			b => dadda_tree_2(1)(36),
			ci => dadda_tree_2(2)(36),
			s => dadda_tree_1(1)(36),
			co => dadda_tree_1(0)(37)
	);
	dadda_tree_1(2)(36) <= dadda_tree_2(3)(36);

	fa_2_0_37: fa
		port map(
			a => dadda_tree_2(0)(37),
			b => dadda_tree_2(1)(37),
			ci => dadda_tree_2(2)(37),
			s => dadda_tree_1(1)(37),
			co => dadda_tree_1(0)(38)
	);
	dadda_tree_1(2)(37) <= dadda_tree_2(3)(37);

	ha_2_0_38: ha
		port map(
			a => dadda_tree_2(0)(38),
			b => dadda_tree_2(1)(38),
			s => dadda_tree_1(1)(38),
			co => dadda_tree_1(0)(39)
	);

	dadda_tree_1(2)(38) <= dadda_tree_2(2)(38);
	dadda_tree_1(0)(39) <= dadda_tree_2(0)(39);
	dadda_tree_1(0)(40) <= dadda_tree_2(0)(40);
	dadda_tree_1(1)(40) <= dadda_tree_2(1)(40);
	dadda_tree_1(0)(41) <= dadda_tree_2(0)(41);
	dadda_tree_1(1)(41) <= dadda_tree_2(1)(41);
	dadda_tree_1(2)(41) <= dadda_tree_2(2)(41);
	dadda_tree_1(0)(42) <= dadda_tree_2(0)(42);
	dadda_tree_1(1)(42) <= dadda_tree_2(1)(42);
	dadda_tree_1(0)(43) <= dadda_tree_2(0)(43);
	dadda_tree_1(1)(43) <= dadda_tree_2(1)(43);
	dadda_tree_1(0)(44) <= dadda_tree_2(0)(44);
	dadda_tree_1(0)(45) <= dadda_tree_2(0)(45);
	dadda_tree_1(1)(45) <= dadda_tree_2(1)(45);
	dadda_tree_1(2)(45) <= dadda_tree_2(2)(45);

	ha_2_0_46: ha
		port map(
			a => dadda_tree_2(0)(46),
			b => dadda_tree_2(1)(46),
			s => dadda_tree_1(0)(46),
			co => dadda_tree_1(0)(47)
	);

	dadda_tree_1(1)(46) <= dadda_tree_2(2)(46);
	dadda_tree_1(2)(46) <= dadda_tree_2(3)(46);

	fa_2_0_47: fa
		port map(
			a => dadda_tree_2(0)(47),
			b => dadda_tree_2(1)(47),
			ci => dadda_tree_2(2)(47),
			s => dadda_tree_1(1)(47),
			co => dadda_tree_1(0)(48)
	);
	dadda_tree_1(2)(47) <= dadda_tree_2(3)(47);

	ha_2_0_48: ha
		port map(
			a => dadda_tree_2(0)(48),
			b => dadda_tree_2(1)(48),
			s => dadda_tree_1(1)(48),
			co => dadda_tree_1(0)(49)
	);

	dadda_tree_1(2)(48) <= dadda_tree_2(2)(48);

	ha_2_0_49: ha
		port map(
			a => dadda_tree_2(0)(49),
			b => dadda_tree_2(1)(49),
			s => dadda_tree_1(1)(49),
			co => dadda_tree_1(0)(50)
	);

	dadda_tree_1(2)(49) <= dadda_tree_2(2)(49);
	dadda_tree_1(0)(50) <= dadda_tree_2(0)(50);
	dadda_tree_1(1)(50) <= dadda_tree_2(1)(50);
	dadda_tree_1(0)(51) <= dadda_tree_2(0)(51);
	dadda_tree_1(0)(52) <= dadda_tree_2(0)(52);
	dadda_tree_1(1)(52) <= dadda_tree_2(1)(52);
	dadda_tree_1(2)(52) <= dadda_tree_2(2)(52);

	ha_2_0_53: ha
		port map(
			a => dadda_tree_2(0)(53),
			b => dadda_tree_2(1)(53),
			s => dadda_tree_1(0)(53),
			co => dadda_tree_1(0)(54)
	);

	dadda_tree_1(1)(53) <= dadda_tree_2(2)(53);
	dadda_tree_1(2)(53) <= dadda_tree_2(3)(53);

	fa_2_0_54: fa
		port map(
			a => dadda_tree_2(0)(54),
			b => dadda_tree_2(1)(54),
			ci => dadda_tree_2(2)(54),
			s => dadda_tree_1(1)(54),
			co => dadda_tree_1(0)(55)
	);
	dadda_tree_1(2)(54) <= dadda_tree_2(3)(54);

	ha_2_0_55: ha
		port map(
			a => dadda_tree_2(0)(55),
			b => dadda_tree_2(1)(55),
			s => dadda_tree_1(1)(55),
			co => dadda_tree_1(0)(56)
	);

	dadda_tree_1(2)(55) <= dadda_tree_2(2)(55);
	dadda_tree_1(0)(56) <= dadda_tree_2(0)(56);
	dadda_tree_1(1)(56) <= dadda_tree_2(1)(56);
	dadda_tree_1(0)(57) <= dadda_tree_2(0)(57);
	dadda_tree_1(0)(58) <= dadda_tree_2(0)(58);
	dadda_tree_1(1)(58) <= dadda_tree_2(1)(58);
	dadda_tree_1(0)(59) <= dadda_tree_2(0)(59);
	dadda_tree_1(1)(59) <= dadda_tree_2(1)(59);
	dadda_tree_1(0)(60) <= dadda_tree_2(0)(60);
	dadda_tree_1(1)(60) <= dadda_tree_2(1)(60);
	dadda_tree_1(0)(61) <= dadda_tree_2(0)(61);
	dadda_tree_1(1)(61) <= dadda_tree_2(1)(61);
	dadda_tree_1(2)(61) <= dadda_tree_2(2)(61);
	dadda_tree_1(0)(62) <= dadda_tree_2(0)(62);
	dadda_tree_1(1)(62) <= dadda_tree_2(1)(62);
	dadda_tree_1(2)(62) <= dadda_tree_2(2)(62);
	dadda_tree_1(0)(63) <= dadda_tree_2(0)(63);
	dadda_tree_1(1)(63) <= dadda_tree_2(1)(63);
	dadda_tree_0(0)(0) <= dadda_tree_1(0)(0);
	dadda_tree_0(1)(0) <= dadda_tree_1(1)(0);
	dadda_tree_0(0)(1) <= dadda_tree_1(0)(1);

	ha_1_0_2: ha
		port map(
			a => dadda_tree_1(0)(2),
			b => dadda_tree_1(1)(2),
			s => dadda_tree_0(0)(2),
			co => dadda_tree_0(0)(3)
	);

	dadda_tree_0(1)(2) <= dadda_tree_1(2)(2);

	ha_1_0_3: ha
		port map(
			a => dadda_tree_1(0)(3),
			b => dadda_tree_1(1)(3),
			s => dadda_tree_0(1)(3),
			co => dadda_tree_0(0)(4)
	);

	dadda_tree_0(0)(4) <= dadda_tree_1(0)(4);
	dadda_tree_0(0)(5) <= dadda_tree_1(0)(5);
	dadda_tree_0(1)(5) <= dadda_tree_1(1)(5);
	dadda_tree_0(0)(6) <= dadda_tree_1(0)(6);
	dadda_tree_0(0)(7) <= dadda_tree_1(0)(7);
	dadda_tree_0(1)(7) <= dadda_tree_1(1)(7);

	ha_1_0_8: ha
		port map(
			a => dadda_tree_1(0)(8),
			b => dadda_tree_1(1)(8),
			s => dadda_tree_0(0)(8),
			co => dadda_tree_0(0)(9)
	);

	dadda_tree_0(1)(8) <= dadda_tree_1(2)(8);
	dadda_tree_0(0)(9) <= dadda_tree_1(0)(9);
	dadda_tree_0(0)(10) <= dadda_tree_1(0)(10);
	dadda_tree_0(0)(11) <= dadda_tree_1(0)(11);
	dadda_tree_0(1)(11) <= dadda_tree_1(1)(11);

	ha_1_0_12: ha
		port map(
			a => dadda_tree_1(0)(12),
			b => dadda_tree_1(1)(12),
			s => dadda_tree_0(0)(12),
			co => dadda_tree_0(0)(13)
	);

	dadda_tree_0(1)(12) <= dadda_tree_1(2)(12);
	dadda_tree_0(0)(13) <= dadda_tree_1(0)(13);
	dadda_tree_0(0)(14) <= dadda_tree_1(0)(14);

	ha_1_0_15: ha
		port map(
			a => dadda_tree_1(0)(15),
			b => dadda_tree_1(1)(15),
			s => dadda_tree_0(0)(15),
			co => dadda_tree_0(0)(16)
	);

	dadda_tree_0(1)(15) <= dadda_tree_1(2)(15);
	dadda_tree_0(0)(16) <= dadda_tree_1(0)(16);
	dadda_tree_0(0)(17) <= dadda_tree_1(0)(17);
	dadda_tree_0(1)(17) <= dadda_tree_1(1)(17);

	ha_1_0_18: ha
		port map(
			a => dadda_tree_1(0)(18),
			b => dadda_tree_1(1)(18),
			s => dadda_tree_0(0)(18),
			co => dadda_tree_0(0)(19)
	);

	dadda_tree_0(1)(18) <= dadda_tree_1(2)(18);
	dadda_tree_0(0)(19) <= dadda_tree_1(0)(19);
	dadda_tree_0(0)(20) <= dadda_tree_1(0)(20);

	ha_1_0_21: ha
		port map(
			a => dadda_tree_1(0)(21),
			b => dadda_tree_1(1)(21),
			s => dadda_tree_0(0)(21),
			co => dadda_tree_0(0)(22)
	);

	dadda_tree_0(1)(21) <= dadda_tree_1(2)(21);
	dadda_tree_0(0)(22) <= dadda_tree_1(0)(22);

	ha_1_0_23: ha
		port map(
			a => dadda_tree_1(0)(23),
			b => dadda_tree_1(1)(23),
			s => dadda_tree_0(0)(23),
			co => dadda_tree_0(0)(24)
	);

	dadda_tree_0(1)(23) <= dadda_tree_1(2)(23);
	dadda_tree_0(0)(24) <= dadda_tree_1(0)(24);
	dadda_tree_0(0)(25) <= dadda_tree_1(0)(25);
	dadda_tree_0(1)(25) <= dadda_tree_1(1)(25);

	ha_1_0_26: ha
		port map(
			a => dadda_tree_1(0)(26),
			b => dadda_tree_1(1)(26),
			s => dadda_tree_0(0)(26),
			co => dadda_tree_0(0)(27)
	);

	dadda_tree_0(1)(26) <= dadda_tree_1(2)(26);
	dadda_tree_0(0)(27) <= dadda_tree_1(0)(27);
	dadda_tree_0(0)(28) <= dadda_tree_1(0)(28);

	ha_1_0_29: ha
		port map(
			a => dadda_tree_1(0)(29),
			b => dadda_tree_1(1)(29),
			s => dadda_tree_0(0)(29),
			co => dadda_tree_0(0)(30)
	);

	dadda_tree_0(1)(29) <= dadda_tree_1(2)(29);
	dadda_tree_0(0)(30) <= dadda_tree_1(0)(30);

	ha_1_0_31: ha
		port map(
			a => dadda_tree_1(0)(31),
			b => dadda_tree_1(1)(31),
			s => dadda_tree_0(0)(31),
			co => dadda_tree_0(0)(32)
	);

	dadda_tree_0(1)(31) <= dadda_tree_1(2)(31);
	dadda_tree_0(0)(32) <= dadda_tree_1(0)(32);
	dadda_tree_0(0)(33) <= dadda_tree_1(0)(33);
	dadda_tree_0(1)(33) <= dadda_tree_1(1)(33);
	dadda_tree_0(0)(34) <= dadda_tree_1(0)(34);
	dadda_tree_0(1)(34) <= dadda_tree_1(1)(34);
	dadda_tree_0(0)(35) <= dadda_tree_1(0)(35);
	dadda_tree_0(1)(35) <= dadda_tree_1(1)(35);
	dadda_tree_0(0)(36) <= dadda_tree_1(0)(36);
	dadda_tree_0(1)(36) <= dadda_tree_1(1)(36);
	dadda_tree_0(0)(37) <= dadda_tree_1(0)(37);
	dadda_tree_0(1)(37) <= dadda_tree_1(1)(37);
	dadda_tree_0(0)(38) <= dadda_tree_1(0)(38);
	dadda_tree_0(1)(38) <= dadda_tree_1(1)(38);
	dadda_tree_0(0)(39) <= dadda_tree_1(0)(39);
	dadda_tree_0(0)(40) <= dadda_tree_1(0)(40);
	dadda_tree_0(1)(40) <= dadda_tree_1(1)(40);

	ha_1_0_41: ha
		port map(
			a => dadda_tree_1(0)(41),
			b => dadda_tree_1(1)(41),
			s => dadda_tree_0(0)(41),
			co => dadda_tree_0(0)(42)
	);

	dadda_tree_0(1)(41) <= dadda_tree_1(2)(41);

	ha_1_0_42: ha
		port map(
			a => dadda_tree_1(0)(42),
			b => dadda_tree_1(1)(42),
			s => dadda_tree_0(1)(42),
			co => dadda_tree_0(0)(43)
	);


	ha_1_0_43: ha
		port map(
			a => dadda_tree_1(0)(43),
			b => dadda_tree_1(1)(43),
			s => dadda_tree_0(1)(43),
			co => dadda_tree_0(0)(44)
	);

	dadda_tree_0(0)(44) <= dadda_tree_1(0)(44);

	ha_1_0_45: ha
		port map(
			a => dadda_tree_1(0)(45),
			b => dadda_tree_1(1)(45),
			s => dadda_tree_0(0)(45),
			co => dadda_tree_0(0)(46)
	);

	dadda_tree_0(1)(45) <= dadda_tree_1(2)(45);
	dadda_tree_0(0)(46) <= dadda_tree_1(0)(46);
	dadda_tree_0(0)(47) <= dadda_tree_1(0)(47);
	dadda_tree_0(1)(47) <= dadda_tree_1(1)(47);
	dadda_tree_0(0)(48) <= dadda_tree_1(0)(48);
	dadda_tree_0(1)(48) <= dadda_tree_1(1)(48);
	dadda_tree_0(0)(49) <= dadda_tree_1(0)(49);
	dadda_tree_0(1)(49) <= dadda_tree_1(1)(49);
	dadda_tree_0(0)(50) <= dadda_tree_1(0)(50);
	dadda_tree_0(1)(50) <= dadda_tree_1(1)(50);
	dadda_tree_0(0)(51) <= dadda_tree_1(0)(51);

	ha_1_0_52: ha
		port map(
			a => dadda_tree_1(0)(52),
			b => dadda_tree_1(1)(52),
			s => dadda_tree_0(0)(52),
			co => dadda_tree_0(0)(53)
	);

	dadda_tree_0(1)(52) <= dadda_tree_1(2)(52);
	dadda_tree_0(0)(53) <= dadda_tree_1(0)(53);
	dadda_tree_0(0)(54) <= dadda_tree_1(0)(54);
	dadda_tree_0(1)(54) <= dadda_tree_1(1)(54);
	dadda_tree_0(0)(55) <= dadda_tree_1(0)(55);
	dadda_tree_0(1)(55) <= dadda_tree_1(1)(55);
	dadda_tree_0(0)(56) <= dadda_tree_1(0)(56);
	dadda_tree_0(1)(56) <= dadda_tree_1(1)(56);
	dadda_tree_0(0)(57) <= dadda_tree_1(0)(57);
	dadda_tree_0(0)(58) <= dadda_tree_1(0)(58);
	dadda_tree_0(1)(58) <= dadda_tree_1(1)(58);
	dadda_tree_0(0)(59) <= dadda_tree_1(0)(59);
	dadda_tree_0(1)(59) <= dadda_tree_1(1)(59);
	dadda_tree_0(0)(60) <= dadda_tree_1(0)(60);
	dadda_tree_0(1)(60) <= dadda_tree_1(1)(60);

	ha_1_0_61: ha
		port map(
			a => dadda_tree_1(0)(61),
			b => dadda_tree_1(1)(61),
			s => dadda_tree_0(0)(61),
			co => dadda_tree_0(0)(62)
	);

	dadda_tree_0(1)(61) <= dadda_tree_1(2)(61);

	fa_1_0_62: fa
		port map(
			a => dadda_tree_1(0)(62),
			b => dadda_tree_1(1)(62),
			ci => dadda_tree_1(2)(62),
			s => dadda_tree_0(1)(62),
			co => dadda_tree_0(0)(63)
	);

	ha_1_0_63: ha
		port map(
			a => dadda_tree_1(0)(63),
			b => dadda_tree_1(1)(63),
			s => dadda_tree_0(1)(63),
			co => open
	);
	dadda_tree_0(1)(1) <= '0';
	dadda_tree_0(1)(2) <= '0';
	dadda_tree_0(1)(4) <= '0';
	dadda_tree_0(1)(6) <= '0';
	dadda_tree_0(1)(8) <= '0';
	dadda_tree_0(1)(9) <= '0';
	dadda_tree_0(1)(10) <= '0';
	dadda_tree_0(1)(12) <= '0';
	dadda_tree_0(1)(13) <= '0';
	dadda_tree_0(1)(14) <= '0';
	dadda_tree_0(1)(15) <= '0';
	dadda_tree_0(1)(16) <= '0';
	dadda_tree_0(1)(18) <= '0';
	dadda_tree_0(1)(19) <= '0';
	dadda_tree_0(1)(20) <= '0';
	dadda_tree_0(1)(21) <= '0';
	dadda_tree_0(1)(22) <= '0';
	dadda_tree_0(1)(23) <= '0';
	dadda_tree_0(1)(24) <= '0';
	dadda_tree_0(1)(26) <= '0';
	dadda_tree_0(1)(27) <= '0';
	dadda_tree_0(1)(28) <= '0';
	dadda_tree_0(1)(29) <= '0';
	dadda_tree_0(1)(30) <= '0';
	dadda_tree_0(1)(31) <= '0';
	dadda_tree_0(1)(32) <= '0';
	dadda_tree_0(1)(39) <= '0';
	dadda_tree_0(1)(41) <= '0';
	dadda_tree_0(1)(44) <= '0';
	dadda_tree_0(1)(45) <= '0';
	dadda_tree_0(1)(46) <= '0';
	dadda_tree_0(1)(51) <= '0';
	dadda_tree_0(1)(52) <= '0';
	dadda_tree_0(1)(53) <= '0';
	dadda_tree_0(1)(57) <= '0';
	dadda_tree_0(1)(61) <= '0';


end architecture structural;